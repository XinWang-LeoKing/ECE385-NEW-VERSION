//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  10-06-2017                               --
//                                                                       --
//    Fall 2017 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 8                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

// This color mapper is for the background

// color_mapper: Decide which color to be output to VGA for each pixel.
module  color_mapper (input [9:0] DrawX, DrawY, // Current pixel coordinates
                      input [11:0] spriteColor, // for background
							 input [7:0] spriteColor_tracer_1, spriteColor_tracer_2, // for tracer
							 input is_tracer_1, is_tracer_2, // current pixel belongs to tracer or not
							 input [23:0] bullet_color,dart_color_center, dart_color_body,
							 input is_healthbar, 
							 input [1:0] chara_id_1, chara_id_2,
							 input [9:0] count_k_1, count_k_2, count_l_1, count_l_2, 
							 input is_energybar,
                      
                      output logic [7:0] VGA_R, VGA_G, VGA_B // VGA RGB output
							 );
    
    logic [7:0] Red, Green, Blue;
    
    // Output colors to VGA
    assign VGA_R = Red;
    assign VGA_G = Green;
    assign VGA_B = Blue;

    // Assign color based on the coordinate
    always_comb
    begin
			if (is_healthbar)
			begin
				Red = 8'h0;
				Green = 8'hff;
				Blue = 8'h0;
			end
			else if (is_energybar)
			begin
				Red = 8'h0;
				Green = 8'h0;
				Blue = 8'hff;
			end
			else if (is_tracer_1&&spriteColor_tracer_1!=0)// draw character 1
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_tracer_1)
8'h0:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'h1:begin Red = 8'h00;Green = 8'h00;Blue = 8'h00;end
8'h2:begin Red = 8'hfa;Green = 8'hce;Blue = 8'ha8;end
8'h3:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha9;end
8'h4:begin Red = 8'hf2;Green = 8'h9d;Blue = 8'h32;end
8'h5:begin Red = 8'hf1;Green = 8'h9e;Blue = 8'h32;end
8'h6:begin Red = 8'hf3;Green = 8'h7e;Blue = 8'h11;end
8'h7:begin Red = 8'hf3;Green = 8'h9e;Blue = 8'h32;end
8'h8:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha8;end
8'h9:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha8;end
8'ha:begin Red = 8'hf2;Green = 8'h9e;Blue = 8'h33;end
8'hb:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha7;end
8'hc:begin Red = 8'h49;Green = 8'h44;Blue = 8'h40;end
8'hd:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hd0;end
8'he:begin Red = 8'hd7;Green = 8'hd1;Blue = 8'hcf;end
8'hf:begin Red = 8'hd7;Green = 8'hd2;Blue = 8'hd0;end
8'h10:begin Red = 8'hd6;Green = 8'hd0;Blue = 8'hce;end
8'h11:begin Red = 8'h47;Green = 8'h42;Blue = 8'h3f;end
8'h12:begin Red = 8'hfb;Green = 8'hcd;Blue = 8'ha7;end
8'h13:begin Red = 8'h87;Green = 8'h62;Blue = 8'h47;end
8'h14:begin Red = 8'h87;Green = 8'h62;Blue = 8'h46;end
8'h15:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hf1;end
8'h16:begin Red = 8'hd6;Green = 8'hcf;Blue = 8'hcd;end
8'h17:begin Red = 8'hd7;Green = 8'hd0;Blue = 8'hce;end
8'h18:begin Red = 8'h55;Green = 8'h39;Blue = 8'h26;end
8'h19:begin Red = 8'h54;Green = 8'h39;Blue = 8'h25;end
8'h1a:begin Red = 8'h86;Green = 8'h61;Blue = 8'h46;end
8'h1b:begin Red = 8'h87;Green = 8'h62;Blue = 8'h45;end
8'h1c:begin Red = 8'h6a;Green = 8'h66;Blue = 8'h62;end
8'h1d:begin Red = 8'h6c;Green = 8'h66;Blue = 8'h64;end
8'h1e:begin Red = 8'hf1;Green = 8'h9d;Blue = 8'h31;end
8'h1f:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hea;end
8'h20:begin Red = 8'hf3;Green = 8'hee;Blue = 8'heb;end
8'h21:begin Red = 8'hf2;Green = 8'hed;Blue = 8'heb;end
8'h22:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hec;end
8'h23:begin Red = 8'h69;Green = 8'h66;Blue = 8'h61;end
8'h24:begin Red = 8'hbc;Green = 8'hb9;Blue = 8'hbb;end
8'h25:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbd;end
8'h26:begin Red = 8'hbb;Green = 8'hba;Blue = 8'hbc;end
8'h27:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbc;end
8'h28:begin Red = 8'hbc;Green = 8'hb8;Blue = 8'hba;end
8'h29:begin Red = 8'h87;Green = 8'h62;Blue = 8'h48;end
8'h2a:begin Red = 8'h55;Green = 8'h39;Blue = 8'h28;end
8'h2b:begin Red = 8'h54;Green = 8'h39;Blue = 8'h26;end
8'h2c:begin Red = 8'h41;Green = 8'h4f;Blue = 8'h61;end
8'h2d:begin Red = 8'h54;Green = 8'h39;Blue = 8'h28;end
8'h2e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h46;end
8'h2f:begin Red = 8'hf3;Green = 8'hed;Blue = 8'heb;end
8'h30:begin Red = 8'hf4;Green = 8'hed;Blue = 8'heb;end
8'h31:begin Red = 8'hf3;Green = 8'hec;Blue = 8'heb;end
8'h32:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbb;end
8'h33:begin Red = 8'h88;Green = 8'h63;Blue = 8'h47;end
8'h34:begin Red = 8'h55;Green = 8'h39;Blue = 8'h27;end
8'h35:begin Red = 8'h56;Green = 8'h39;Blue = 8'h28;end
8'h36:begin Red = 8'h53;Green = 8'h39;Blue = 8'h25;end
8'h37:begin Red = 8'h55;Green = 8'h38;Blue = 8'h27;end
8'h38:begin Red = 8'h86;Green = 8'h61;Blue = 8'h45;end
8'h39:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd8;end
8'h3a:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd7;end
8'h3b:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd8;end
8'h3c:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd9;end
8'h3d:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd8;end
8'h3e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h48;end
8'h3f:begin Red = 8'h88;Green = 8'h63;Blue = 8'h48;end
8'h40:begin Red = 8'h88;Green = 8'h62;Blue = 8'h47;end
8'h41:begin Red = 8'h6b;Green = 8'h66;Blue = 8'h63;end
8'h42:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd9;end
8'h43:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hd9;end
8'h44:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hda;end
8'h45:begin Red = 8'h86;Green = 8'h61;Blue = 8'h47;end
8'h46:begin Red = 8'h86;Green = 8'h60;Blue = 8'h45;end
8'h47:begin Red = 8'hda;Green = 8'hd8;Blue = 8'hd9;end
8'h48:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd9;end
8'h49:begin Red = 8'h42;Green = 8'h4f;Blue = 8'h61;end
8'h4a:begin Red = 8'h87;Green = 8'h61;Blue = 8'h46;end
8'h4b:begin Red = 8'h87;Green = 8'h61;Blue = 8'h47;end
8'h4c:begin Red = 8'h41;Green = 8'h50;Blue = 8'h62;end
8'h4d:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h44;end
8'h4e:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1c;end
8'h4f:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h22;end
8'h50:begin Red = 8'hf6;Green = 8'h9b;Blue = 8'h11;end
8'h51:begin Red = 8'hf8;Green = 8'h9d;Blue = 8'h14;end
8'h52:begin Red = 8'hf6;Green = 8'h7e;Blue = 8'h18;end
8'h53:begin Red = 8'hf7;Green = 8'h80;Blue = 8'h18;end
8'h54:begin Red = 8'hf3;Green = 8'heb;Blue = 8'he9;end
8'h55:begin Red = 8'hf3;Green = 8'hee;Blue = 8'hec;end
8'h56:begin Red = 8'hf2;Green = 8'heb;Blue = 8'hea;end
8'h57:begin Red = 8'hf3;Green = 8'heb;Blue = 8'hea;end
8'h58:begin Red = 8'hf3;Green = 8'hed;Blue = 8'hea;end
8'h59:begin Red = 8'hd9;Green = 8'hd5;Blue = 8'hd8;end
8'h5a:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1a;end
8'h5b:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h1a;end
8'h5c:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h19;end
8'h5d:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h16;end
8'h5e:begin Red = 8'hfa;Green = 8'hc2;Blue = 8'h1a;end
8'h5f:begin Red = 8'h41;Green = 8'h4e;Blue = 8'h60;end
8'h60:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h17;end
8'h61:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h43;end
8'h62:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h17;end
8'h63:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h43;end
8'h64:begin Red = 8'h42;Green = 8'h51;Blue = 8'h63;end
8'h65:begin Red = 8'hf9;Green = 8'hc2;Blue = 8'h19;end
8'h66:begin Red = 8'hb5;Green = 8'h9a;Blue = 8'h44;end
8'h67:begin Red = 8'h40;Green = 8'h4e;Blue = 8'h60;end
8'h68:begin Red = 8'hb5;Green = 8'h99;Blue = 8'h43;end
8'h69:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h1a;end
8'h6a:begin Red = 8'he2;Green = 8'ha2;Blue = 8'h22;end
8'h6b:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h44;end
8'h6c:begin Red = 8'hf7;Green = 8'h9c;Blue = 8'h14;end
8'h6d:begin Red = 8'hf7;Green = 8'h9b;Blue = 8'h14;end
8'h6e:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h42;end
8'h6f:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h43;end
8'h70:begin Red = 8'hb3;Green = 8'h99;Blue = 8'h43;end
8'h71:begin Red = 8'hf6;Green = 8'h9c;Blue = 8'h14;end
8'h72:begin Red = 8'hf7;Green = 8'h9d;Blue = 8'h14;end
8'h73:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h19;end
8'h74:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h22;end
8'h75:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h20;end
8'h76:begin Red = 8'he0;Green = 8'ha1;Blue = 8'h22;end
8'h77:begin Red = 8'he1;Green = 8'ha3;Blue = 8'h21;end
8'h78:begin Red = 8'hf6;Green = 8'h7d;Blue = 8'h16;end
8'h79:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h23;end
8'h7a:begin Red = 8'hf8;Green = 8'h9e;Blue = 8'h14;end
8'h7b:begin Red = 8'he1;Green = 8'ha1;Blue = 8'h20;end
8'h7c:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h21;end
8'h7d:begin Red = 8'he2;Green = 8'ha4;Blue = 8'h22;end
8'h7e:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h1b;end
8'h7f:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h1a;end
8'h80:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h18;end
8'h81:begin Red = 8'h71;Green = 8'h92;Blue = 8'hff;end
8'h82:begin Red = 8'hfc;Green = 8'hea;Blue = 8'hff;end
8'h83:begin Red = 8'hfd;Green = 8'hea;Blue = 8'hff;end
8'h84:begin Red = 8'hf8;Green = 8'hd5;Blue = 8'hff;end
8'h85:begin Red = 8'hf7;Green = 8'hd6;Blue = 8'hff;end
8'h86:begin Red = 8'hf8;Green = 8'hc8;Blue = 8'hff;end
8'h87:begin Red = 8'hf8;Green = 8'hd6;Blue = 8'hff;end
8'h88:begin Red = 8'h9a;Green = 8'haf;Blue = 8'hff;end
8'h89:begin Red = 8'he8;Green = 8'hc7;Blue = 8'hff;end
8'h8a:begin Red = 8'he9;Green = 8'heb;Blue = 8'hff;end
8'h8b:begin Red = 8'he9;Green = 8'hec;Blue = 8'hff;end
8'h8c:begin Red = 8'he8;Green = 8'heb;Blue = 8'hff;end
8'h8d:begin Red = 8'h99;Green = 8'hae;Blue = 8'hff;end
8'h8e:begin Red = 8'hbc;Green = 8'hbc;Blue = 8'hff;end
8'h8f:begin Red = 8'he8;Green = 8'hc8;Blue = 8'hff;end
8'h90:begin Red = 8'he8;Green = 8'hea;Blue = 8'hff;end
8'h91:begin Red = 8'ha0;Green = 8'haa;Blue = 8'hff;end
8'h92:begin Red = 8'hbc;Green = 8'hbb;Blue = 8'hff;end
8'h93:begin Red = 8'hac;Green = 8'hbe;Blue = 8'hff;end
8'h94:begin Red = 8'had;Green = 8'hbe;Blue = 8'hff;end
8'h95:begin Red = 8'hf7;Green = 8'hd5;Blue = 8'hff;end
8'h96:begin Red = 8'hf8;Green = 8'hf7;Blue = 8'hff;end
8'h97:begin Red = 8'hf8;Green = 8'hf8;Blue = 8'hff;end
8'h98:begin Red = 8'hab;Green = 8'hbe;Blue = 8'hff;end
8'h99:begin Red = 8'hda;Green = 8'he1;Blue = 8'hff;end
8'h9a:begin Red = 8'hda;Green = 8'he2;Blue = 8'hff;end
8'h9b:begin Red = 8'hd9;Green = 8'he2;Blue = 8'hff;end
8'h9c:begin Red = 8'h95;Green = 8'hb4;Blue = 8'hff;end
8'h9d:begin Red = 8'hf9;Green = 8'hf7;Blue = 8'hff;end
8'h9e:begin Red = 8'hbd;Green = 8'hbc;Blue = 8'hff;end
8'h9f:begin Red = 8'ha1;Green = 8'haa;Blue = 8'hff;end
8'ha0:begin Red = 8'h9f;Green = 8'haa;Blue = 8'hff;end
8'ha1:begin Red = 8'hea;Green = 8'hee;Blue = 8'hff;end
8'ha2:begin Red = 8'hea;Green = 8'hed;Blue = 8'hff;end
8'ha3:begin Red = 8'h96;Green = 8'hb4;Blue = 8'hff;end
8'ha4:begin Red = 8'hd5;Green = 8'hd4;Blue = 8'hff;end
8'ha5:begin Red = 8'hfc;Green = 8'he4;Blue = 8'hff;end
8'ha6:begin Red = 8'hee;Green = 8'hd7;Blue = 8'hff;end
8'ha7:begin Red = 8'hfa;Green = 8'hd4;Blue = 8'hff;end
8'ha8:begin Red = 8'hfb;Green = 8'hd5;Blue = 8'hff;end
8'ha9:begin Red = 8'hfa;Green = 8'hc8;Blue = 8'hff;end
8'haa:begin Red = 8'hfb;Green = 8'hc9;Blue = 8'hff;end
8'hab:begin Red = 8'hf8;Green = 8'hf6;Blue = 8'hff;end
8'hac:begin Red = 8'hfc;Green = 8'he5;Blue = 8'hff;end
8'had:begin Red = 8'h95;Green = 8'hb3;Blue = 8'hff;end
8'hae:begin Red = 8'hd5;Green = 8'hd3;Blue = 8'hff;end
8'haf:begin Red = 8'h96;Green = 8'hb5;Blue = 8'hff;end
8'hb0:begin Red = 8'hd6;Green = 8'hd4;Blue = 8'hff;end
8'hb1:begin Red = 8'hd6;Green = 8'hd3;Blue = 8'hff;end
8'hb2:begin Red = 8'hef;Green = 8'hd7;Blue = 8'hff;end
8'hb3:begin Red = 8'hfb;Green = 8'hd4;Blue = 8'hff;end
8'hb4:begin Red = 8'hfa;Green = 8'hd5;Blue = 8'hff;end
8'hb5:begin Red = 8'hfb;Green = 8'hc8;Blue = 8'hff;end
8'hb6:begin Red = 8'hef;Green = 8'hd8;Blue = 8'hff;end
8'hb7:begin Red = 8'hee;Green = 8'hd8;Blue = 8'hff;end
8'hb8:begin Red = 8'hfa;Green = 8'hc7;Blue = 8'hff;end
8'hb9:begin Red = 8'hfb;Green = 8'hd6;Blue = 8'hff;end
endcase
			end
			else if (is_tracer_2&&spriteColor_tracer_2!=0) // draw character 2
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_tracer_2)
8'h0:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'h1:begin Red = 8'h00;Green = 8'h00;Blue = 8'h00;end
8'h2:begin Red = 8'hfa;Green = 8'hce;Blue = 8'ha8;end
8'h3:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha9;end
8'h4:begin Red = 8'hf2;Green = 8'h9d;Blue = 8'h32;end
8'h5:begin Red = 8'hf1;Green = 8'h9e;Blue = 8'h32;end
8'h6:begin Red = 8'hf3;Green = 8'h7e;Blue = 8'h11;end
8'h7:begin Red = 8'hf3;Green = 8'h9e;Blue = 8'h32;end
8'h8:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha8;end
8'h9:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha8;end
8'ha:begin Red = 8'hf2;Green = 8'h9e;Blue = 8'h33;end
8'hb:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha7;end
8'hc:begin Red = 8'h49;Green = 8'h44;Blue = 8'h40;end
8'hd:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hd0;end
8'he:begin Red = 8'hd7;Green = 8'hd1;Blue = 8'hcf;end
8'hf:begin Red = 8'hd7;Green = 8'hd2;Blue = 8'hd0;end
8'h10:begin Red = 8'hd6;Green = 8'hd0;Blue = 8'hce;end
8'h11:begin Red = 8'h47;Green = 8'h42;Blue = 8'h3f;end
8'h12:begin Red = 8'hfb;Green = 8'hcd;Blue = 8'ha7;end
8'h13:begin Red = 8'h87;Green = 8'h62;Blue = 8'h47;end
8'h14:begin Red = 8'h87;Green = 8'h62;Blue = 8'h46;end
8'h15:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hf1;end
8'h16:begin Red = 8'hd6;Green = 8'hcf;Blue = 8'hcd;end
8'h17:begin Red = 8'hd7;Green = 8'hd0;Blue = 8'hce;end
8'h18:begin Red = 8'h55;Green = 8'h39;Blue = 8'h26;end
8'h19:begin Red = 8'h54;Green = 8'h39;Blue = 8'h25;end
8'h1a:begin Red = 8'h86;Green = 8'h61;Blue = 8'h46;end
8'h1b:begin Red = 8'h87;Green = 8'h62;Blue = 8'h45;end
8'h1c:begin Red = 8'h6a;Green = 8'h66;Blue = 8'h62;end
8'h1d:begin Red = 8'h6c;Green = 8'h66;Blue = 8'h64;end
8'h1e:begin Red = 8'hf1;Green = 8'h9d;Blue = 8'h31;end
8'h1f:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hea;end
8'h20:begin Red = 8'hf3;Green = 8'hee;Blue = 8'heb;end
8'h21:begin Red = 8'hf2;Green = 8'hed;Blue = 8'heb;end
8'h22:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hec;end
8'h23:begin Red = 8'h69;Green = 8'h66;Blue = 8'h61;end
8'h24:begin Red = 8'hbc;Green = 8'hb9;Blue = 8'hbb;end
8'h25:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbd;end
8'h26:begin Red = 8'hbb;Green = 8'hba;Blue = 8'hbc;end
8'h27:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbc;end
8'h28:begin Red = 8'hbc;Green = 8'hb8;Blue = 8'hba;end
8'h29:begin Red = 8'h87;Green = 8'h62;Blue = 8'h48;end
8'h2a:begin Red = 8'h55;Green = 8'h39;Blue = 8'h28;end
8'h2b:begin Red = 8'h54;Green = 8'h39;Blue = 8'h26;end
8'h2c:begin Red = 8'h41;Green = 8'h4f;Blue = 8'h61;end
8'h2d:begin Red = 8'h54;Green = 8'h39;Blue = 8'h28;end
8'h2e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h46;end
8'h2f:begin Red = 8'hf3;Green = 8'hed;Blue = 8'heb;end
8'h30:begin Red = 8'hf4;Green = 8'hed;Blue = 8'heb;end
8'h31:begin Red = 8'hf3;Green = 8'hec;Blue = 8'heb;end
8'h32:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbb;end
8'h33:begin Red = 8'h88;Green = 8'h63;Blue = 8'h47;end
8'h34:begin Red = 8'h55;Green = 8'h39;Blue = 8'h27;end
8'h35:begin Red = 8'h56;Green = 8'h39;Blue = 8'h28;end
8'h36:begin Red = 8'h53;Green = 8'h39;Blue = 8'h25;end
8'h37:begin Red = 8'h55;Green = 8'h38;Blue = 8'h27;end
8'h38:begin Red = 8'h86;Green = 8'h61;Blue = 8'h45;end
8'h39:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd8;end
8'h3a:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd7;end
8'h3b:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd8;end
8'h3c:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd9;end
8'h3d:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd8;end
8'h3e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h48;end
8'h3f:begin Red = 8'h88;Green = 8'h63;Blue = 8'h48;end
8'h40:begin Red = 8'h88;Green = 8'h62;Blue = 8'h47;end
8'h41:begin Red = 8'h6b;Green = 8'h66;Blue = 8'h63;end
8'h42:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd9;end
8'h43:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hd9;end
8'h44:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hda;end
8'h45:begin Red = 8'h86;Green = 8'h61;Blue = 8'h47;end
8'h46:begin Red = 8'h86;Green = 8'h60;Blue = 8'h45;end
8'h47:begin Red = 8'hda;Green = 8'hd8;Blue = 8'hd9;end
8'h48:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd9;end
8'h49:begin Red = 8'h42;Green = 8'h4f;Blue = 8'h61;end
8'h4a:begin Red = 8'h87;Green = 8'h61;Blue = 8'h46;end
8'h4b:begin Red = 8'h87;Green = 8'h61;Blue = 8'h47;end
8'h4c:begin Red = 8'h41;Green = 8'h50;Blue = 8'h62;end
8'h4d:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h44;end
8'h4e:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1c;end
8'h4f:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h22;end
8'h50:begin Red = 8'hf6;Green = 8'h9b;Blue = 8'h11;end
8'h51:begin Red = 8'hf8;Green = 8'h9d;Blue = 8'h14;end
8'h52:begin Red = 8'hf6;Green = 8'h7e;Blue = 8'h18;end
8'h53:begin Red = 8'hf7;Green = 8'h80;Blue = 8'h18;end
8'h54:begin Red = 8'hf3;Green = 8'heb;Blue = 8'he9;end
8'h55:begin Red = 8'hf3;Green = 8'hee;Blue = 8'hec;end
8'h56:begin Red = 8'hf2;Green = 8'heb;Blue = 8'hea;end
8'h57:begin Red = 8'hf3;Green = 8'heb;Blue = 8'hea;end
8'h58:begin Red = 8'hf3;Green = 8'hed;Blue = 8'hea;end
8'h59:begin Red = 8'hd9;Green = 8'hd5;Blue = 8'hd8;end
8'h5a:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1a;end
8'h5b:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h1a;end
8'h5c:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h19;end
8'h5d:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h16;end
8'h5e:begin Red = 8'hfa;Green = 8'hc2;Blue = 8'h1a;end
8'h5f:begin Red = 8'h41;Green = 8'h4e;Blue = 8'h60;end
8'h60:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h17;end
8'h61:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h43;end
8'h62:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h17;end
8'h63:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h43;end
8'h64:begin Red = 8'h42;Green = 8'h51;Blue = 8'h63;end
8'h65:begin Red = 8'hf9;Green = 8'hc2;Blue = 8'h19;end
8'h66:begin Red = 8'hb5;Green = 8'h9a;Blue = 8'h44;end
8'h67:begin Red = 8'h40;Green = 8'h4e;Blue = 8'h60;end
8'h68:begin Red = 8'hb5;Green = 8'h99;Blue = 8'h43;end
8'h69:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h1a;end
8'h6a:begin Red = 8'he2;Green = 8'ha2;Blue = 8'h22;end
8'h6b:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h44;end
8'h6c:begin Red = 8'hf7;Green = 8'h9c;Blue = 8'h14;end
8'h6d:begin Red = 8'hf7;Green = 8'h9b;Blue = 8'h14;end
8'h6e:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h42;end
8'h6f:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h43;end
8'h70:begin Red = 8'hb3;Green = 8'h99;Blue = 8'h43;end
8'h71:begin Red = 8'hf6;Green = 8'h9c;Blue = 8'h14;end
8'h72:begin Red = 8'hf7;Green = 8'h9d;Blue = 8'h14;end
8'h73:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h19;end
8'h74:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h22;end
8'h75:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h20;end
8'h76:begin Red = 8'he0;Green = 8'ha1;Blue = 8'h22;end
8'h77:begin Red = 8'he1;Green = 8'ha3;Blue = 8'h21;end
8'h78:begin Red = 8'hf6;Green = 8'h7d;Blue = 8'h16;end
8'h79:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h23;end
8'h7a:begin Red = 8'hf8;Green = 8'h9e;Blue = 8'h14;end
8'h7b:begin Red = 8'he1;Green = 8'ha1;Blue = 8'h20;end
8'h7c:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h21;end
8'h7d:begin Red = 8'he2;Green = 8'ha4;Blue = 8'h22;end
8'h7e:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h1b;end
8'h7f:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h1a;end
8'h80:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h18;end
8'h81:begin Red = 8'h71;Green = 8'h92;Blue = 8'hff;end
8'h82:begin Red = 8'hfc;Green = 8'hea;Blue = 8'hff;end
8'h83:begin Red = 8'hfd;Green = 8'hea;Blue = 8'hff;end
8'h84:begin Red = 8'hf8;Green = 8'hd5;Blue = 8'hff;end
8'h85:begin Red = 8'hf7;Green = 8'hd6;Blue = 8'hff;end
8'h86:begin Red = 8'hf8;Green = 8'hc8;Blue = 8'hff;end
8'h87:begin Red = 8'hf8;Green = 8'hd6;Blue = 8'hff;end
8'h88:begin Red = 8'h9a;Green = 8'haf;Blue = 8'hff;end
8'h89:begin Red = 8'he8;Green = 8'hc7;Blue = 8'hff;end
8'h8a:begin Red = 8'he9;Green = 8'heb;Blue = 8'hff;end
8'h8b:begin Red = 8'he9;Green = 8'hec;Blue = 8'hff;end
8'h8c:begin Red = 8'he8;Green = 8'heb;Blue = 8'hff;end
8'h8d:begin Red = 8'h99;Green = 8'hae;Blue = 8'hff;end
8'h8e:begin Red = 8'hbc;Green = 8'hbc;Blue = 8'hff;end
8'h8f:begin Red = 8'he8;Green = 8'hc8;Blue = 8'hff;end
8'h90:begin Red = 8'he8;Green = 8'hea;Blue = 8'hff;end
8'h91:begin Red = 8'ha0;Green = 8'haa;Blue = 8'hff;end
8'h92:begin Red = 8'hbc;Green = 8'hbb;Blue = 8'hff;end
8'h93:begin Red = 8'hac;Green = 8'hbe;Blue = 8'hff;end
8'h94:begin Red = 8'had;Green = 8'hbe;Blue = 8'hff;end
8'h95:begin Red = 8'hf7;Green = 8'hd5;Blue = 8'hff;end
8'h96:begin Red = 8'hf8;Green = 8'hf7;Blue = 8'hff;end
8'h97:begin Red = 8'hf8;Green = 8'hf8;Blue = 8'hff;end
8'h98:begin Red = 8'hab;Green = 8'hbe;Blue = 8'hff;end
8'h99:begin Red = 8'hda;Green = 8'he1;Blue = 8'hff;end
8'h9a:begin Red = 8'hda;Green = 8'he2;Blue = 8'hff;end
8'h9b:begin Red = 8'hd9;Green = 8'he2;Blue = 8'hff;end
8'h9c:begin Red = 8'h95;Green = 8'hb4;Blue = 8'hff;end
8'h9d:begin Red = 8'hf9;Green = 8'hf7;Blue = 8'hff;end
8'h9e:begin Red = 8'hbd;Green = 8'hbc;Blue = 8'hff;end
8'h9f:begin Red = 8'ha1;Green = 8'haa;Blue = 8'hff;end
8'ha0:begin Red = 8'h9f;Green = 8'haa;Blue = 8'hff;end
8'ha1:begin Red = 8'hea;Green = 8'hee;Blue = 8'hff;end
8'ha2:begin Red = 8'hea;Green = 8'hed;Blue = 8'hff;end
8'ha3:begin Red = 8'h96;Green = 8'hb4;Blue = 8'hff;end
8'ha4:begin Red = 8'hd5;Green = 8'hd4;Blue = 8'hff;end
8'ha5:begin Red = 8'hfc;Green = 8'he4;Blue = 8'hff;end
8'ha6:begin Red = 8'hee;Green = 8'hd7;Blue = 8'hff;end
8'ha7:begin Red = 8'hfa;Green = 8'hd4;Blue = 8'hff;end
8'ha8:begin Red = 8'hfb;Green = 8'hd5;Blue = 8'hff;end
8'ha9:begin Red = 8'hfa;Green = 8'hc8;Blue = 8'hff;end
8'haa:begin Red = 8'hfb;Green = 8'hc9;Blue = 8'hff;end
8'hab:begin Red = 8'hf8;Green = 8'hf6;Blue = 8'hff;end
8'hac:begin Red = 8'hfc;Green = 8'he5;Blue = 8'hff;end
8'had:begin Red = 8'h95;Green = 8'hb3;Blue = 8'hff;end
8'hae:begin Red = 8'hd5;Green = 8'hd3;Blue = 8'hff;end
8'haf:begin Red = 8'h96;Green = 8'hb5;Blue = 8'hff;end
8'hb0:begin Red = 8'hd6;Green = 8'hd4;Blue = 8'hff;end
8'hb1:begin Red = 8'hd6;Green = 8'hd3;Blue = 8'hff;end
8'hb2:begin Red = 8'hef;Green = 8'hd7;Blue = 8'hff;end
8'hb3:begin Red = 8'hfb;Green = 8'hd4;Blue = 8'hff;end
8'hb4:begin Red = 8'hfa;Green = 8'hd5;Blue = 8'hff;end
8'hb5:begin Red = 8'hfb;Green = 8'hc8;Blue = 8'hff;end
8'hb6:begin Red = 8'hef;Green = 8'hd8;Blue = 8'hff;end
8'hb7:begin Red = 8'hee;Green = 8'hd8;Blue = 8'hff;end
8'hb8:begin Red = 8'hfa;Green = 8'hc7;Blue = 8'hff;end
8'hb9:begin Red = 8'hfb;Green = 8'hd6;Blue = 8'hff;end
endcase
			end
			else if (bullet_color!=24'h000000) begin
					Red = bullet_color[23:16];
					Green = bullet_color[15:8];
					Blue = bullet_color[7:0];
			end
			/*else if (dart_color_body==24'hffff00)begin
					Red = dart_color_body[23:16];
					Green = dart_color_body[15:8];
					Blue = dart_color_body[7:0];
			end
			else if (dart_color_center==24'hffffff)begin
					Red = dart_color_center[23:16];
					Green = dart_color_center[15:8];
					Blue = dart_color_center[7:0];
			end*/
			//else if ((bullet_state==2'b01||bullet_state==2'b10)&&bullet_x==DrawX&&bullet_y==DrawY)
			/*else if(bullet_x>=DrawX-1'b1&&bullet_x<=DrawX+1'b1&&bullet_y>=DrawY-1'b1&&bullet_y<=DrawY+1'b1)
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'h00;	
			end*/
			else // draw background
			begin
				  Red   = 8'hff;
				  Green = 8'h00;
				  Blue  = 8'h00;
				  /*case(spriteColor)
12'h0:    begin Red = 8'h3c;    Green = 8'h58;    Blue = 8'h5f;
end 12'h1:    begin Red = 8'h3f;    Green = 8'h5c;    Blue = 8'h64;
end 12'h2:    begin Red = 8'h29;    Green = 8'h44;    Blue = 8'h4b;
end 12'h3:    begin Red = 8'h2f;    Green = 8'h4a;    Blue = 8'h51;
end 12'h4:    begin Red = 8'h89;    Green = 8'hf5;    Blue = 8'hfe;
end 12'h5:    begin Red = 8'h81;    Green = 8'hdc;    Blue = 8'hf6;
end 12'h6:    begin Red = 8'h73;    Green = 8'hdb;    Blue = 8'he3;
end 12'h7:    begin Red = 8'h71;    Green = 8'hc0;    Blue = 8'hdd;
end 12'h8:    begin Red = 8'h73;    Green = 8'hc1;    Blue = 8'hd6;
end 12'h9:    begin Red = 8'h75;    Green = 8'hd1;    Blue = 8'he7;
end 12'ha:    begin Red = 8'h7a;    Green = 8'hd0;    Blue = 8'he8;
end 12'hb:    begin Red = 8'h79;    Green = 8'hda;    Blue = 8'hf9;
end 12'hc:    begin Red = 8'h60;    Green = 8'h7d;    Blue = 8'h77;
end 12'hd:    begin Red = 8'h65;    Green = 8'h82;    Blue = 8'h87;
end 12'he:    begin Red = 8'h52;    Green = 8'h80;    Blue = 8'h75;
end 12'hf:    begin Red = 8'h5e;    Green = 8'h7c;    Blue = 8'h7d;
end 12'h10:    begin Red = 8'h32;    Green = 8'h4f;    Blue = 8'h57;
end 12'h11:    begin Red = 8'h36;    Green = 8'h54;    Blue = 8'h5d;
end 12'h12:    begin Red = 8'h26;    Green = 8'h37;    Blue = 8'h3f;
end 12'h13:    begin Red = 8'h2d;    Green = 8'h40;    Blue = 8'h46;
end 12'h14:    begin Red = 8'h28;    Green = 8'h2a;    Blue = 8'h39;
end 12'h15:    begin Red = 8'h71;    Green = 8'hc3;    Blue = 8'hd0;
end 12'h16:    begin Red = 8'h6d;    Green = 8'hc6;    Blue = 8'hd5;
end 12'h17:    begin Red = 8'h5f;    Green = 8'h81;    Blue = 8'h81;
end 12'h18:    begin Red = 8'h55;    Green = 8'h71;    Blue = 8'h73;
end 12'h19:    begin Red = 8'h24;    Green = 8'h32;    Blue = 8'h32;
end 12'h1a:    begin Red = 8'h26;    Green = 8'h28;    Blue = 8'h34;
end 12'h1b:    begin Red = 8'h19;    Green = 8'h2c;    Blue = 8'h30;
end 12'h1c:    begin Red = 8'h79;    Green = 8'hbb;    Blue = 8'hdd;
end 12'h1d:    begin Red = 8'h5b;    Green = 8'h5e;    Blue = 8'h53;
end 12'h1e:    begin Red = 8'h5c;    Green = 8'h6a;    Blue = 8'h6a;
end 12'h1f:    begin Red = 8'h64;    Green = 8'h7d;    Blue = 8'h83;
end 12'h20:    begin Red = 8'h5a;    Green = 8'h81;    Blue = 8'h7b;
end 12'h21:    begin Red = 8'h2b;    Green = 8'h4d;    Blue = 8'h4c;
end 12'h22:    begin Red = 8'h2e;    Green = 8'h4a;    Blue = 8'h57;
end 12'h23:    begin Red = 8'h36;    Green = 8'h47;    Blue = 8'h56;
end 12'h24:    begin Red = 8'h79;    Green = 8'hd4;    Blue = 8'hed;
end 12'h25:    begin Red = 8'h6b;    Green = 8'hc3;    Blue = 8'hce;
end 12'h26:    begin Red = 8'h71;    Green = 8'hba;    Blue = 8'hd9;
end 12'h27:    begin Red = 8'h5d;    Green = 8'h79;    Blue = 8'h83;
end 12'h28:    begin Red = 8'h62;    Green = 8'h78;    Blue = 8'h85;
end 12'h29:    begin Red = 8'h3b;    Green = 8'h59;    Blue = 8'h5a;
end 12'h2a:    begin Red = 8'h2d;    Green = 8'h3d;    Blue = 8'h3c;
end 12'h2b:    begin Red = 8'h36;    Green = 8'h4b;    Blue = 8'h4b;
end 12'h2c:    begin Red = 8'h22;    Green = 8'h4a;    Blue = 8'h48;
end 12'h2d:    begin Red = 8'h31;    Green = 8'h42;    Blue = 8'h51;
end 12'h2e:    begin Red = 8'h6b;    Green = 8'hc0;    Blue = 8'hd3;
end 12'h2f:    begin Red = 8'h61;    Green = 8'h71;    Blue = 8'h70;
end 12'h30:    begin Red = 8'h8f;    Green = 8'haf;    Blue = 8'h85;
end 12'h31:    begin Red = 8'h8b;    Green = 8'hac;    Blue = 8'h80;
end 12'h32:    begin Red = 8'h39;    Green = 8'h54;    Blue = 8'h64;
end 12'h33:    begin Red = 8'h41;    Green = 8'h62;    Blue = 8'h6a;
end 12'h34:    begin Red = 8'h7a;    Green = 8'hdc;    Blue = 8'hf2;
end 12'h35:    begin Red = 8'h76;    Green = 8'hbf;    Blue = 8'hc9;
end 12'h36:    begin Red = 8'h80;    Green = 8'ha0;    Blue = 8'h7a;
end 12'h37:    begin Red = 8'h83;    Green = 8'ha2;    Blue = 8'h7f;
end 12'h38:    begin Red = 8'h23;    Green = 8'h3f;    Blue = 8'h41;
end 12'h39:    begin Red = 8'h2b;    Green = 8'h34;    Blue = 8'h3c;
end 12'h3a:    begin Red = 8'h1e;    Green = 8'h31;    Blue = 8'h2d;
end 12'h3b:    begin Red = 8'h1d;    Green = 8'h17;    Blue = 8'h23;
end 12'h3c:    begin Red = 8'h60;    Green = 8'h61;    Blue = 8'h5b;
end 12'h3d:    begin Red = 8'h57;    Green = 8'h6b;    Blue = 8'h68;
end 12'h3e:    begin Red = 8'h5f;    Green = 8'h77;    Blue = 8'h7a;
end 12'h3f:    begin Red = 8'h89;    Green = 8'haa;    Blue = 8'h78;
end 12'h40:    begin Red = 8'h62;    Green = 8'h77;    Blue = 8'h57;
end 12'h41:    begin Red = 8'h22;    Green = 8'h35;    Blue = 8'h3a;
end 12'h42:    begin Red = 8'h29;    Green = 8'h51;    Blue = 8'h52;
end 12'h43:    begin Red = 8'h21;    Green = 8'h30;    Blue = 8'h42;
end 12'h44:    begin Red = 8'h6b;    Green = 8'h75;    Blue = 8'h7e;
end 12'h45:    begin Red = 8'h5a;    Green = 8'h77;    Blue = 8'h7c;
end 12'h46:    begin Red = 8'h57;    Green = 8'h72;    Blue = 8'h82;
end 12'h47:    begin Red = 8'h84;    Green = 8'ha8;    Blue = 8'h74;
end 12'h48:    begin Red = 8'h84;    Green = 8'ha3;    Blue = 8'h74;
end 12'h49:    begin Red = 8'h5a;    Green = 8'h72;    Blue = 8'h57;
end 12'h4a:    begin Red = 8'h65;    Green = 8'h79;    Blue = 8'h5f;
end 12'h4b:    begin Red = 8'h21;    Green = 8'h3a;    Blue = 8'h3e;
end 12'h4c:    begin Red = 8'h2f;    Green = 8'h4c;    Blue = 8'h47;
end 12'h4d:    begin Red = 8'h59;    Green = 8'h76;    Blue = 8'h76;
end 12'h4e:    begin Red = 8'h89;    Green = 8'hab;    Blue = 8'h89;
end 12'h4f:    begin Red = 8'h8f;    Green = 8'hab;    Blue = 8'h8b;
end 12'h50:    begin Red = 8'h60;    Green = 8'h79;    Blue = 8'h5e;
end 12'h51:    begin Red = 8'h47;    Green = 8'h5f;    Blue = 8'h63;
end 12'h52:    begin Red = 8'h1b;    Green = 8'h38;    Blue = 8'h3b;
end 12'h53:    begin Red = 8'h81;    Green = 8'h9d;    Blue = 8'h80;
end 12'h54:    begin Red = 8'h86;    Green = 8'ha3;    Blue = 8'h86;
end 12'h55:    begin Red = 8'h8b;    Green = 8'ha5;    Blue = 8'h85;
end 12'h56:    begin Red = 8'h96;    Green = 8'hae;    Blue = 8'h8f;
end 12'h57:    begin Red = 8'h63;    Green = 8'h7e;    Blue = 8'h56;
end 12'h58:    begin Red = 8'h44;    Green = 8'h56;    Blue = 8'h61;
end 12'h59:    begin Red = 8'hd3;    Green = 8'hcf;    Blue = 8'hbe;
end 12'h5a:    begin Red = 8'hbc;    Green = 8'hb8;    Blue = 8'ha7;
end 12'h5b:    begin Red = 8'hbc;    Green = 8'hb3;    Blue = 8'ha4;
end 12'h5c:    begin Red = 8'hc9;    Green = 8'hc0;    Blue = 8'hb1;
end 12'h5d:    begin Red = 8'hc3;    Green = 8'hbc;    Blue = 8'hab;
end 12'h5e:    begin Red = 8'h3e;    Green = 8'h55;    Blue = 8'h65;
end 12'h5f:    begin Red = 8'hb9;    Green = 8'hb8;    Blue = 8'hac;
end 12'h60:    begin Red = 8'ha6;    Green = 8'ha5;    Blue = 8'h99;
end 12'h61:    begin Red = 8'h34;    Green = 8'h4d;    Blue = 8'h51;
end 12'h62:    begin Red = 8'hb4;    Green = 8'hb8;    Blue = 8'hb2;
end 12'h63:    begin Red = 8'h57;    Green = 8'h72;    Blue = 8'h7d;
end 12'h64:    begin Red = 8'h57;    Green = 8'h70;    Blue = 8'h52;
end 12'h65:    begin Red = 8'h5f;    Green = 8'h7f;    Blue = 8'h86;
end 12'h66:    begin Red = 8'h33;    Green = 8'h51;    Blue = 8'h64;
end 12'h67:    begin Red = 8'h3b;    Green = 8'h56;    Blue = 8'h6a;
end 12'h68:    begin Red = 8'h1c;    Green = 8'h46;    Blue = 8'h50;
end 12'h69:    begin Red = 8'h23;    Green = 8'h48;    Blue = 8'h60;
end 12'h6a:    begin Red = 8'h24;    Green = 8'h44;    Blue = 8'h51;
end 12'h6b:    begin Red = 8'hac;    Green = 8'hb2;    Blue = 8'ha8;
end 12'h6c:    begin Red = 8'ha8;    Green = 8'hb5;    Blue = 8'ha1;
end 12'h6d:    begin Red = 8'h6a;    Green = 8'h88;    Blue = 8'h88;
end 12'h6e:    begin Red = 8'h5d;    Green = 8'h7c;    Blue = 8'h70;
end 12'h6f:    begin Red = 8'h62;    Green = 8'h74;    Blue = 8'h5d;
end 12'h70:    begin Red = 8'h71;    Green = 8'h80;    Blue = 8'h52;
end 12'h71:    begin Red = 8'h2a;    Green = 8'h57;    Blue = 8'h54;
end 12'h72:    begin Red = 8'h91;    Green = 8'h6f;    Blue = 8'h4f;
end 12'h73:    begin Red = 8'ha9;    Green = 8'ha7;    Blue = 8'ha0;
end 12'h74:    begin Red = 8'ha2;    Green = 8'ha6;    Blue = 8'ha0;
end 12'h75:    begin Red = 8'h87;    Green = 8'h66;    Blue = 8'h3d;
end 12'h76:    begin Red = 8'h8d;    Green = 8'h99;    Blue = 8'h8e;
end 12'h77:    begin Red = 8'h8f;    Green = 8'h87;    Blue = 8'h72;
end 12'h78:    begin Red = 8'ha2;    Green = 8'ha1;    Blue = 8'h94;
end 12'h79:    begin Red = 8'h81;    Green = 8'h9d;    Blue = 8'h89;
end 12'h7a:    begin Red = 8'h85;    Green = 8'ha4;    Blue = 8'h79;
end 12'h7b:    begin Red = 8'h59;    Green = 8'h6e;    Blue = 8'h61;
end 12'h7c:    begin Red = 8'h60;    Green = 8'h78;    Blue = 8'h64;
end 12'h7d:    begin Red = 8'h30;    Green = 8'h48;    Blue = 8'h4c;
end 12'h7e:    begin Red = 8'ha5;    Green = 8'h7e;    Blue = 8'h4e;
end 12'h7f:    begin Red = 8'ha7;    Green = 8'h83;    Blue = 8'h58;
end 12'h80:    begin Red = 8'h96;    Green = 8'h71;    Blue = 8'h4c;
end 12'h81:    begin Red = 8'haf;    Green = 8'ha6;    Blue = 8'ha0;
end 12'h82:    begin Red = 8'haa;    Green = 8'haa;    Blue = 8'h9a;
end 12'h83:    begin Red = 8'hbf;    Green = 8'hbe;    Blue = 8'hb1;
end 12'h84:    begin Red = 8'h7e;    Green = 8'h63;    Blue = 8'h47;
end 12'h85:    begin Red = 8'h8c;    Green = 8'h72;    Blue = 8'h49;
end 12'h86:    begin Red = 8'h94;    Green = 8'h8d;    Blue = 8'h7f;
end 12'h87:    begin Red = 8'h87;    Green = 8'h86;    Blue = 8'h7a;
end 12'h88:    begin Red = 8'h32;    Green = 8'h4a;    Blue = 8'h5d;
end 12'h89:    begin Red = 8'hae;    Green = 8'h7f;    Blue = 8'h5a;
end 12'h8a:    begin Red = 8'h82;    Green = 8'h63;    Blue = 8'h40;
end 12'h8b:    begin Red = 8'h8d;    Green = 8'h73;    Blue = 8'h54;
end 12'h8c:    begin Red = 8'h8d;    Green = 8'h8f;    Blue = 8'h7c;
end 12'h8d:    begin Red = 8'h89;    Green = 8'h84;    Blue = 8'h69;
end 12'h8e:    begin Red = 8'hae;    Green = 8'ha2;    Blue = 8'h99;
end 12'h8f:    begin Red = 8'hc2;    Green = 8'h84;    Blue = 8'h57;
end 12'h90:    begin Red = 8'h93;    Green = 8'h6b;    Blue = 8'h3f;
end 12'h91:    begin Red = 8'h90;    Green = 8'h6a;    Blue = 8'h4e;
end 12'h92:    begin Red = 8'h9e;    Green = 8'ha7;    Blue = 8'h99;
end 12'h93:    begin Red = 8'h10;    Green = 8'h3e;    Blue = 8'h4b;
end 12'h94:    begin Red = 8'hb6;    Green = 8'h93;    Blue = 8'h6b;
end 12'h95:    begin Red = 8'hbd;    Green = 8'h96;    Blue = 8'h6d;
end 12'h96:    begin Red = 8'h52;    Green = 8'h7d;    Blue = 8'h7c;
end 12'h97:    begin Red = 8'h64;    Green = 8'h78;    Blue = 8'h77;
end 12'h98:    begin Red = 8'h4e;    Green = 8'h6b;    Blue = 8'h6b;
end 12'h99:    begin Red = 8'h55;    Green = 8'h6c;    Blue = 8'h74;
end 12'h9a:    begin Red = 8'h98;    Green = 8'hba;    Blue = 8'h73;
end 12'h9b:    begin Red = 8'h6f;    Green = 8'h81;    Blue = 8'h5f;
end 12'h9c:    begin Red = 8'h74;    Green = 8'h86;    Blue = 8'h57;
end 12'h9d:    begin Red = 8'ha8;    Green = 8'h7d;    Blue = 8'h56;
end 12'h9e:    begin Red = 8'h92;    Green = 8'h91;    Blue = 8'h84;
end 12'h9f:    begin Red = 8'ha2;    Green = 8'ha2;    Blue = 8'h8f;
end 12'ha0:    begin Red = 8'h77;    Green = 8'h76;    Blue = 8'h68;
end 12'ha1:    begin Red = 8'h15;    Green = 8'h39;    Blue = 8'h43;
end 12'ha2:    begin Red = 8'haa;    Green = 8'h8c;    Blue = 8'h6a;
end 12'ha3:    begin Red = 8'haa;    Green = 8'h90;    Blue = 8'h6f;
end 12'ha4:    begin Red = 8'h9a;    Green = 8'h99;    Blue = 8'h8c;
end 12'ha5:    begin Red = 8'h97;    Green = 8'h96;    Blue = 8'h87;
end 12'ha6:    begin Red = 8'h9b;    Green = 8'h6d;    Blue = 8'h43;
end 12'ha7:    begin Red = 8'h7f;    Green = 8'h7c;    Blue = 8'h6e;
end 12'ha8:    begin Red = 8'h90;    Green = 8'h78;    Blue = 8'h54;
end 12'ha9:    begin Red = 8'ha1;    Green = 8'h99;    Blue = 8'h79;
end 12'haa:    begin Red = 8'hb1;    Green = 8'h8f;    Blue = 8'h64;
end 12'hab:    begin Red = 8'hab;    Green = 8'h90;    Blue = 8'h75;
end 12'hac:    begin Red = 8'ha5;    Green = 8'h90;    Blue = 8'h75;
end 12'had:    begin Red = 8'h8b;    Green = 8'h7c;    Blue = 8'h60;
end 12'hae:    begin Red = 8'h69;    Green = 8'h83;    Blue = 8'h58;
end 12'haf:    begin Red = 8'h90;    Green = 8'h6d;    Blue = 8'h49;
end 12'hb0:    begin Red = 8'h14;    Green = 8'h39;    Blue = 8'h4b;
end 12'hb1:    begin Red = 8'h06;    Green = 8'h34;    Blue = 8'h4f;
end 12'hb2:    begin Red = 8'h91;    Green = 8'h7e;    Blue = 8'h64;
end 12'hb3:    begin Red = 8'haf;    Green = 8'h95;    Blue = 8'h73;
end 12'hb4:    begin Red = 8'haa;    Green = 8'h91;    Blue = 8'h69;
end 12'hb5:    begin Red = 8'hae;    Green = 8'h97;    Blue = 8'h6e;
end 12'hb6:    begin Red = 8'h4c;    Green = 8'h75;    Blue = 8'h80;
end 12'hb7:    begin Red = 8'h54;    Green = 8'h71;    Blue = 8'h67;
end 12'hb8:    begin Red = 8'h4c;    Green = 8'h66;    Blue = 8'h6b;
end 12'hb9:    begin Red = 8'h30;    Green = 8'h4f;    Blue = 8'h5c;
end 12'hba:    begin Red = 8'h90;    Green = 8'h64;    Blue = 8'h39;
end 12'hbb:    begin Red = 8'h8d;    Green = 8'h77;    Blue = 8'h5a;
end 12'hbc:    begin Red = 8'haf;    Green = 8'h8f;    Blue = 8'h70;
end 12'hbd:    begin Red = 8'h4d;    Green = 8'h67;    Blue = 8'h70;
end 12'hbe:    begin Red = 8'h68;    Green = 8'h7e;    Blue = 8'h62;
end 12'hbf:    begin Red = 8'h92;    Green = 8'h79;    Blue = 8'h5f;
end 12'hc0:    begin Red = 8'h59;    Green = 8'h72;    Blue = 8'h88;
end 12'hc1:    begin Red = 8'h39;    Green = 8'h5c;    Blue = 8'h4d;
end 12'hc2:    begin Red = 8'h3d;    Green = 8'h5c;    Blue = 8'h69;
end 12'hc3:    begin Red = 8'hf3;    Green = 8'hea;    Blue = 8'haf;
end 12'hc4:    begin Red = 8'hdb;    Green = 8'hd4;    Blue = 8'ha9;
end 12'hc5:    begin Red = 8'hd9;    Green = 8'hd9;    Blue = 8'had;
end 12'hc6:    begin Red = 8'h88;    Green = 8'h90;    Blue = 8'h7c;
end 12'hc7:    begin Red = 8'h8e;    Green = 8'h96;    Blue = 8'h80;
end 12'hc8:    begin Red = 8'h77;    Green = 8'h7e;    Blue = 8'h6c;
end 12'hc9:    begin Red = 8'h74;    Green = 8'h85;    Blue = 8'h72;
end 12'hca:    begin Red = 8'h7a;    Green = 8'h85;    Blue = 8'h74;
end 12'hcb:    begin Red = 8'ha6;    Green = 8'ha7;    Blue = 8'h8f;
end 12'hcc:    begin Red = 8'h7d;    Green = 8'h7f;    Blue = 8'h68;
end 12'hcd:    begin Red = 8'h6c;    Green = 8'h79;    Blue = 8'h5e;
end 12'hce:    begin Red = 8'h72;    Green = 8'h7c;    Blue = 8'h69;
end 12'hcf:    begin Red = 8'h73;    Green = 8'h7c;    Blue = 8'h62;
end 12'hd0:    begin Red = 8'h6c;    Green = 8'h6b;    Blue = 8'h5f;
end 12'hd1:    begin Red = 8'h6f;    Green = 8'h61;    Blue = 8'h56;
end 12'hd2:    begin Red = 8'h5f;    Green = 8'h62;    Blue = 8'h48;
end 12'hd3:    begin Red = 8'h85;    Green = 8'h84;    Blue = 8'h75;
end 12'hd4:    begin Red = 8'h1d;    Green = 8'h44;    Blue = 8'h4b;
end 12'hd5:    begin Red = 8'h01;    Green = 8'h2c;    Blue = 8'h3d;
end 12'hd6:    begin Red = 8'h08;    Green = 8'h29;    Blue = 8'h38;
end 12'hd7:    begin Red = 8'h4d;    Green = 8'h6d;    Blue = 8'h73;
end 12'hd8:    begin Red = 8'h35;    Green = 8'h65;    Blue = 8'h70;
end 12'hd9:    begin Red = 8'h38;    Green = 8'h68;    Blue = 8'h76;
end 12'hda:    begin Red = 8'h3e;    Green = 8'h67;    Blue = 8'h70;
end 12'hdb:    begin Red = 8'h44;    Green = 8'h67;    Blue = 8'h72;
end 12'hdc:    begin Red = 8'h53;    Green = 8'h6c;    Blue = 8'h80;
end 12'hdd:    begin Red = 8'h5e;    Green = 8'h7e;    Blue = 8'h51;
end 12'hde:    begin Red = 8'he2;    Green = 8'hd4;    Blue = 8'ha1;
end 12'hdf:    begin Red = 8'hc0;    Green = 8'hbe;    Blue = 8'ha1;
end 12'he0:    begin Red = 8'hb9;    Green = 8'hb9;    Blue = 8'h91;
end 12'he1:    begin Red = 8'h92;    Green = 8'h90;    Blue = 8'h72;
end 12'he2:    begin Red = 8'h7a;    Green = 8'h84;    Blue = 8'h62;
end 12'he3:    begin Red = 8'h82;    Green = 8'h7c;    Blue = 8'h66;
end 12'he4:    begin Red = 8'h7e;    Green = 8'h72;    Blue = 8'h5c;
end 12'he5:    begin Red = 8'h79;    Green = 8'h77;    Blue = 8'h61;
end 12'he6:    begin Red = 8'h89;    Green = 8'h74;    Blue = 8'h6a;
end 12'he7:    begin Red = 8'h67;    Green = 8'h68;    Blue = 8'h59;
end 12'he8:    begin Red = 8'h67;    Green = 8'h66;    Blue = 8'h4d;
end 12'he9:    begin Red = 8'hae;    Green = 8'hac;    Blue = 8'h9f;
end 12'hea:    begin Red = 8'h35;    Green = 8'h46;    Blue = 8'h47;
end 12'heb:    begin Red = 8'hf0;    Green = 8'hd3;    Blue = 8'ha4;
end 12'hec:    begin Red = 8'hb2;    Green = 8'h92;    Blue = 8'h78;
end 12'hed:    begin Red = 8'hb9;    Green = 8'h95;    Blue = 8'h66;
end 12'hee:    begin Red = 8'h5a;    Green = 8'h7c;    Blue = 8'h75;
end 12'hef:    begin Red = 8'hfa;    Green = 8'he7;    Blue = 8'haf;
end 12'hf0:    begin Red = 8'hed;    Green = 8'hd3;    Blue = 8'ha9;
end 12'hf1:    begin Red = 8'h88;    Green = 8'h9e;    Blue = 8'h7c;
end 12'hf2:    begin Red = 8'h88;    Green = 8'ha4;    Blue = 8'h7e;
end 12'hf3:    begin Red = 8'h7e;    Green = 8'ha0;    Blue = 8'h72;
end 12'hf4:    begin Red = 8'h87;    Green = 8'h9d;    Blue = 8'h83;
end 12'hf5:    begin Red = 8'h37;    Green = 8'h5e;    Blue = 8'h54;
end 12'hf6:    begin Red = 8'hd8;    Green = 8'hd2;    Blue = 8'ha2;
end 12'hf7:    begin Red = 8'h85;    Green = 8'h83;    Blue = 8'h6e;
end 12'hf8:    begin Red = 8'hb5;    Green = 8'hb3;    Blue = 8'ha5;
end 12'hf9:    begin Red = 8'h79;    Green = 8'h78;    Blue = 8'h5c;
end 12'hfa:    begin Red = 8'h6e;    Green = 8'h6b;    Blue = 8'h5a;
end 12'hfb:    begin Red = 8'h68;    Green = 8'h65;    Blue = 8'h54;
end 12'hfc:    begin Red = 8'h38;    Green = 8'h49;    Blue = 8'h6c;
end 12'hfd:    begin Red = 8'h8f;    Green = 8'ha2;    Blue = 8'h2a;
end 12'hfe:    begin Red = 8'h8d;    Green = 8'h9d;    Blue = 8'h24;
end 12'hff:    begin Red = 8'hfe;    Green = 8'hfc;    Blue = 8'hc8;
end 12'h100:    begin Red = 8'hff;    Green = 8'hf4;    Blue = 8'hb8;
end 12'h101:    begin Red = 8'hff;    Green = 8'hef;    Blue = 8'hc5;
end 12'h102:    begin Red = 8'hef;    Green = 8'hd8;    Blue = 8'ha7;
end 12'h103:    begin Red = 8'hf6;    Green = 8'hcd;    Blue = 8'h91;
end 12'h104:    begin Red = 8'hf4;    Green = 8'hce;    Blue = 8'h9b;
end 12'h105:    begin Red = 8'ha0;    Green = 8'h95;    Blue = 8'h6a;
end 12'h106:    begin Red = 8'h8c;    Green = 8'h71;    Blue = 8'h4e;
end 12'h107:    begin Red = 8'h58;    Green = 8'h3f;    Blue = 8'h23;
end 12'h108:    begin Red = 8'h5f;    Green = 8'h49;    Blue = 8'h2d;
end 12'h109:    begin Red = 8'h5d;    Green = 8'h45;    Blue = 8'h26;
end 12'h10a:    begin Red = 8'ha7;    Green = 8'h89;    Blue = 8'h72;
end 12'h10b:    begin Red = 8'hec;    Green = 8'hbe;    Blue = 8'h8c;
end 12'h10c:    begin Red = 8'hf2;    Green = 8'hf0;    Blue = 8'hb8;
end 12'h10d:    begin Red = 8'hff;    Green = 8'he7;    Blue = 8'hb0;
end 12'h10e:    begin Red = 8'hff;    Green = 8'hd0;    Blue = 8'ha4;
end 12'h10f:    begin Red = 8'hea;    Green = 8'hd3;    Blue = 8'hb2;
end 12'h110:    begin Red = 8'hff;    Green = 8'hde;    Blue = 8'hab;
end 12'h111:    begin Red = 8'h7a;    Green = 8'h91;    Blue = 8'h71;
end 12'h112:    begin Red = 8'hfc;    Green = 8'hf3;    Blue = 8'hee;
end 12'h113:    begin Red = 8'hf8;    Green = 8'hed;    Blue = 8'hec;
end 12'h114:    begin Red = 8'hff;    Green = 8'hf8;    Blue = 8'hf7;
end 12'h115:    begin Red = 8'h70;    Green = 8'h92;    Blue = 8'h6c;
end 12'h116:    begin Red = 8'h3c;    Green = 8'h59;    Blue = 8'h55;
end 12'h117:    begin Red = 8'h27;    Green = 8'h4f;    Blue = 8'h6c;
end 12'h118:    begin Red = 8'h80;    Green = 8'h8e;    Blue = 8'h35;
end 12'h119:    begin Red = 8'h7c;    Green = 8'h8f;    Blue = 8'h30;
end 12'h11a:    begin Red = 8'hff;    Green = 8'hf1;    Blue = 8'hc0;
end 12'h11b:    begin Red = 8'hf5;    Green = 8'hd0;    Blue = 8'ha4;
end 12'h11c:    begin Red = 8'hed;    Green = 8'hd3;    Blue = 8'h92;
end 12'h11d:    begin Red = 8'hce;    Green = 8'hb3;    Blue = 8'h88;
end 12'h11e:    begin Red = 8'h66;    Green = 8'h4f;    Blue = 8'h37;
end 12'h11f:    begin Red = 8'h6d;    Green = 8'h58;    Blue = 8'h3f;
end 12'h120:    begin Red = 8'hcf;    Green = 8'hb5;    Blue = 8'h82;
end 12'h121:    begin Red = 8'hf6;    Green = 8'hde;    Blue = 8'hb3;
end 12'h122:    begin Red = 8'he6;    Green = 8'hd8;    Blue = 8'hae;
end 12'h123:    begin Red = 8'h92;    Green = 8'h9c;    Blue = 8'h81;
end 12'h124:    begin Red = 8'h63;    Green = 8'h97;    Blue = 8'h62;
end 12'h125:    begin Red = 8'hed;    Green = 8'he1;    Blue = 8'hdd;
end 12'h126:    begin Red = 8'he6;    Green = 8'he1;    Blue = 8'hd7;
end 12'h127:    begin Red = 8'he1;    Green = 8'hdf;    Blue = 8'hda;
end 12'h128:    begin Red = 8'he8;    Green = 8'he6;    Blue = 8'hdd;
end 12'h129:    begin Red = 8'hfe;    Green = 8'heb;    Blue = 8'hf0;
end 12'h12a:    begin Red = 8'hfe;    Green = 8'hed;    Blue = 8'he8;
end 12'h12b:    begin Red = 8'he1;    Green = 8'hde;    Blue = 8'hd5;
end 12'h12c:    begin Red = 8'h6c;    Green = 8'h90;    Blue = 8'h67;
end 12'h12d:    begin Red = 8'h5d;    Green = 8'h7b;    Blue = 8'h59;
end 12'h12e:    begin Red = 8'h63;    Green = 8'h7b;    Blue = 8'h28;
end 12'h12f:    begin Red = 8'h71;    Green = 8'h7e;    Blue = 8'h27;
end 12'h130:    begin Red = 8'h68;    Green = 8'h76;    Blue = 8'h30;
end 12'h131:    begin Red = 8'h66;    Green = 8'h76;    Blue = 8'h26;
end 12'h132:    begin Red = 8'h4d;    Green = 8'h58;    Blue = 8'h1a;
end 12'h133:    begin Red = 8'h3f;    Green = 8'h53;    Blue = 8'h18;
end 12'h134:    begin Red = 8'h7f;    Green = 8'h93;    Blue = 8'h28;
end 12'h135:    begin Red = 8'hfc;    Green = 8'hdf;    Blue = 8'hb0;
end 12'h136:    begin Red = 8'hf5;    Green = 8'hda;    Blue = 8'had;
end 12'h137:    begin Red = 8'hf5;    Green = 8'hd6;    Blue = 8'ha8;
end 12'h138:    begin Red = 8'hff;    Green = 8'he7;    Blue = 8'hbb;
end 12'h139:    begin Red = 8'hc3;    Green = 8'hab;    Blue = 8'h7a;
end 12'h13a:    begin Red = 8'hb8;    Green = 8'h9d;    Blue = 8'h73;
end 12'h13b:    begin Red = 8'hd4;    Green = 8'hb7;    Blue = 8'h89;
end 12'h13c:    begin Red = 8'h97;    Green = 8'h7d;    Blue = 8'h5d;
end 12'h13d:    begin Red = 8'h70;    Green = 8'h57;    Blue = 8'h3a;
end 12'h13e:    begin Red = 8'ha2;    Green = 8'h8b;    Blue = 8'h6a;
end 12'h13f:    begin Red = 8'hd3;    Green = 8'hbc;    Blue = 8'h8c;
end 12'h140:    begin Red = 8'ha5;    Green = 8'h8b;    Blue = 8'h5e;
end 12'h141:    begin Red = 8'hb3;    Green = 8'h9a;    Blue = 8'h6e;
end 12'h142:    begin Red = 8'hef;    Green = 8'hd3;    Blue = 8'h9f;
end 12'h143:    begin Red = 8'he6;    Green = 8'he0;    Blue = 8'hdc;
end 12'h144:    begin Red = 8'he3;    Green = 8'he1;    Blue = 8'he3;
end 12'h145:    begin Red = 8'he5;    Green = 8'hd9;    Blue = 8'hd2;
end 12'h146:    begin Red = 8'hdd;    Green = 8'hd9;    Blue = 8'hd9;
end 12'h147:    begin Red = 8'hfa;    Green = 8'hf0;    Blue = 8'hf3;
end 12'h148:    begin Red = 8'h7f;    Green = 8'h9a;    Blue = 8'h79;
end 12'h149:    begin Red = 8'h67;    Green = 8'h74;    Blue = 8'h63;
end 12'h14a:    begin Red = 8'h3e;    Green = 8'h54;    Blue = 8'h58;
end 12'h14b:    begin Red = 8'hc6;    Green = 8'hc5;    Blue = 8'h98;
end 12'h14c:    begin Red = 8'h33;    Green = 8'h58;    Blue = 8'h6a;
end 12'h14d:    begin Red = 8'h2b;    Green = 8'h4f;    Blue = 8'h76;
end 12'h14e:    begin Red = 8'h2f;    Green = 8'h53;    Blue = 8'h6a;
end 12'h14f:    begin Red = 8'h32;    Green = 8'h51;    Blue = 8'h74;
end 12'h150:    begin Red = 8'h79;    Green = 8'h87;    Blue = 8'h28;
end 12'h151:    begin Red = 8'h71;    Green = 8'h7d;    Blue = 8'h36;
end 12'h152:    begin Red = 8'h66;    Green = 8'h72;    Blue = 8'h2b;
end 12'h153:    begin Red = 8'h48;    Green = 8'h50;    Blue = 8'h1b;
end 12'h154:    begin Red = 8'h3a;    Green = 8'h47;    Blue = 8'h14;
end 12'h155:    begin Red = 8'h88;    Green = 8'h98;    Blue = 8'h21;
end 12'h156:    begin Red = 8'h8c;    Green = 8'h9d;    Blue = 8'h2a;
end 12'h157:    begin Red = 8'hfa;    Green = 8'he4;    Blue = 8'hb7;
end 12'h158:    begin Red = 8'hdc;    Green = 8'hbd;    Blue = 8'h90;
end 12'h159:    begin Red = 8'h85;    Green = 8'h6b;    Blue = 8'h4a;
end 12'h15a:    begin Red = 8'h65;    Green = 8'h4f;    Blue = 8'h31;
end 12'h15b:    begin Red = 8'hb9;    Green = 8'ha1;    Blue = 8'h78;
end 12'h15c:    begin Red = 8'h83;    Green = 8'h6a;    Blue = 8'h50;
end 12'h15d:    begin Red = 8'hd5;    Green = 8'hbd;    Blue = 8'h91;
end 12'h15e:    begin Red = 8'ha6;    Green = 8'h8a;    Blue = 8'h64;
end 12'h15f:    begin Red = 8'h81;    Green = 8'h6a;    Blue = 8'h44;
end 12'h160:    begin Red = 8'hea;    Green = 8'hd2;    Blue = 8'h9f;
end 12'h161:    begin Red = 8'h67;    Green = 8'h96;    Blue = 8'h74;
end 12'h162:    begin Red = 8'h6e;    Green = 8'h8d;    Blue = 8'h5f;
end 12'h163:    begin Red = 8'he9;    Green = 8'he1;    Blue = 8'he3;
end 12'h164:    begin Red = 8'hff;    Green = 8'hf3;    Blue = 8'hf5;
end 12'h165:    begin Red = 8'hf7;    Green = 8'hf8;    Blue = 8'hf2;
end 12'h166:    begin Red = 8'h67;    Green = 8'h6d;    Blue = 8'h59;
end 12'h167:    begin Red = 8'h62;    Green = 8'h6e;    Blue = 8'h5a;
end 12'h168:    begin Red = 8'h70;    Green = 8'h95;    Blue = 8'h64;
end 12'h169:    begin Red = 8'h52;    Green = 8'h6f;    Blue = 8'h49;
end 12'h16a:    begin Red = 8'h45;    Green = 8'h61;    Blue = 8'h41;
end 12'h16b:    begin Red = 8'h5e;    Green = 8'h77;    Blue = 8'h52;
end 12'h16c:    begin Red = 8'h58;    Green = 8'h64;    Blue = 8'h50;
end 12'h16d:    begin Red = 8'h4a;    Green = 8'h63;    Blue = 8'h45;
end 12'h16e:    begin Red = 8'h52;    Green = 8'h68;    Blue = 8'h4c;
end 12'h16f:    begin Red = 8'h45;    Green = 8'h67;    Blue = 8'h51;
end 12'h170:    begin Red = 8'h4b;    Green = 8'h68;    Blue = 8'h45;
end 12'h171:    begin Red = 8'h38;    Green = 8'h4d;    Blue = 8'h60;
end 12'h172:    begin Red = 8'h19;    Green = 8'h3e;    Blue = 8'h46;
end 12'h173:    begin Red = 8'h1a;    Green = 8'h38;    Blue = 8'h4b;
end 12'h174:    begin Red = 8'h92;    Green = 8'h8f;    Blue = 8'h79;
end 12'h175:    begin Red = 8'h4d;    Green = 8'h5a;    Blue = 8'h1f;
end 12'h176:    begin Red = 8'h44;    Green = 8'h56;    Blue = 8'h5a;
end 12'h177:    begin Red = 8'h53;    Green = 8'h5a;    Blue = 8'h1f;
end 12'h178:    begin Red = 8'h67;    Green = 8'h7c;    Blue = 8'h32;
end 12'h179:    begin Red = 8'h3f;    Green = 8'h5d;    Blue = 8'h6e;
end 12'h17a:    begin Red = 8'hf4;    Green = 8'he0;    Blue = 8'hac;
end 12'h17b:    begin Red = 8'h75;    Green = 8'h5d;    Blue = 8'h3a;
end 12'h17c:    begin Red = 8'hc0;    Green = 8'ha0;    Blue = 8'h7a;
end 12'h17d:    begin Red = 8'h6b;    Green = 8'h57;    Blue = 8'h35;
end 12'h17e:    begin Red = 8'hc6;    Green = 8'ha7;    Blue = 8'h82;
end 12'h17f:    begin Red = 8'h60;    Green = 8'h91;    Blue = 8'h70;
end 12'h180:    begin Red = 8'h61;    Green = 8'h7e;    Blue = 8'h62;
end 12'h181:    begin Red = 8'hd5;    Green = 8'hd2;    Blue = 8'hc9;
end 12'h182:    begin Red = 8'hcf;    Green = 8'hcc;    Blue = 8'hc5;
end 12'h183:    begin Red = 8'hf7;    Green = 8'he4;    Blue = 8'hea;
end 12'h184:    begin Red = 8'hd2;    Green = 8'hd6;    Blue = 8'hc3;
end 12'h185:    begin Red = 8'hd9;    Green = 8'hd9;    Blue = 8'hc7;
end 12'h186:    begin Red = 8'hc7;    Green = 8'hcb;    Blue = 8'hbc;
end 12'h187:    begin Red = 8'hd5;    Green = 8'hd0;    Blue = 8'hd4;
end 12'h188:    begin Red = 8'hf4;    Green = 8'hf4;    Blue = 8'he8;
end 12'h189:    begin Red = 8'hd4;    Green = 8'hcd;    Blue = 8'h9f;
end 12'h18a:    begin Red = 8'hc1;    Green = 8'hbf;    Blue = 8'h98;
end 12'h18b:    begin Red = 8'h6b;    Green = 8'h7b;    Blue = 8'h2b;
end 12'h18c:    begin Red = 8'h48;    Green = 8'h59;    Blue = 8'h1f;
end 12'h18d:    begin Red = 8'h52;    Green = 8'h5c;    Blue = 8'h18;
end 12'h18e:    begin Red = 8'h6c;    Green = 8'h7c;    Blue = 8'h34;
end 12'h18f:    begin Red = 8'h2e;    Green = 8'h4d;    Blue = 8'h62;
end 12'h190:    begin Red = 8'h40;    Green = 8'h50;    Blue = 8'h60;
end 12'h191:    begin Red = 8'hc9;    Green = 8'hb4;    Blue = 8'h90;
end 12'h192:    begin Red = 8'h8f;    Green = 8'h78;    Blue = 8'h4f;
end 12'h193:    begin Red = 8'h7a;    Green = 8'h62;    Blue = 8'h41;
end 12'h194:    begin Red = 8'hdc;    Green = 8'hd8;    Blue = 8'hd4;
end 12'h195:    begin Red = 8'hde;    Green = 8'hd9;    Blue = 8'hcf;
end 12'h196:    begin Red = 8'he6;    Green = 8'hdb;    Blue = 8'hd8;
end 12'h197:    begin Red = 8'hc6;    Green = 8'hc6;    Blue = 8'hc0;
end 12'h198:    begin Red = 8'hcc;    Green = 8'hd1;    Blue = 8'hc4;
end 12'h199:    begin Red = 8'hee;    Green = 8'hec;    Blue = 8'heb;
end 12'h19a:    begin Red = 8'h66;    Green = 8'h76;    Blue = 8'h69;
end 12'h19b:    begin Red = 8'hcf;    Green = 8'hca;    Blue = 8'hbe;
end 12'h19c:    begin Red = 8'hcc;    Green = 8'hd0;    Blue = 8'hbf;
end 12'h19d:    begin Red = 8'hce;    Green = 8'hd2;    Blue = 8'hc9;
end 12'h19e:    begin Red = 8'h0b;    Green = 8'h21;    Blue = 8'h2c;
end 12'h19f:    begin Red = 8'h34;    Green = 8'h41;    Blue = 8'h4a;
end 12'h1a0:    begin Red = 8'h4a;    Green = 8'h4e;    Blue = 8'h14;
end 12'h1a1:    begin Red = 8'h4d;    Green = 8'h54;    Blue = 8'h23;
end 12'h1a2:    begin Red = 8'h2b;    Green = 8'h4b;    Blue = 8'h67;
end 12'h1a3:    begin Red = 8'h36;    Green = 8'h5a;    Blue = 8'h5e;
end 12'h1a4:    begin Red = 8'hc4;    Green = 8'hb0;    Blue = 8'h95;
end 12'h1a5:    begin Red = 8'hff;    Green = 8'he5;    Blue = 8'hb6;
end 12'h1a6:    begin Red = 8'h93;    Green = 8'h72;    Blue = 8'h57;
end 12'h1a7:    begin Red = 8'hb5;    Green = 8'h9c;    Blue = 8'h78;
end 12'h1a8:    begin Red = 8'hf8;    Green = 8'heb;    Blue = 8'hf1;
end 12'h1a9:    begin Red = 8'hdc;    Green = 8'hdf;    Blue = 8'hdc;
end 12'h1aa:    begin Red = 8'hce;    Green = 8'hcb;    Blue = 8'hcb;
end 12'h1ab:    begin Red = 8'hf2;    Green = 8'he2;    Blue = 8'hef;
end 12'h1ac:    begin Red = 8'hd8;    Green = 8'hcc;    Blue = 8'hc6;
end 12'h1ad:    begin Red = 8'h8a;    Green = 8'h87;    Blue = 8'h70;
end 12'h1ae:    begin Red = 8'h7c;    Green = 8'h79;    Blue = 8'h67;
end 12'h1af:    begin Red = 8'h02;    Green = 8'hd3;    Blue = 8'hf9;
end 12'h1b0:    begin Red = 8'h03;    Green = 8'h13;    Blue = 8'h2c;
end 12'h1b1:    begin Red = 8'h34;    Green = 8'h3a;    Blue = 8'h19;
end 12'h1b2:    begin Red = 8'h2a;    Green = 8'h31;    Blue = 8'h19;
end 12'h1b3:    begin Red = 8'h4a;    Green = 8'h58;    Blue = 8'h13;
end 12'h1b4:    begin Red = 8'h85;    Green = 8'h9b;    Blue = 8'h39;
end 12'h1b5:    begin Red = 8'h43;    Green = 8'h46;    Blue = 8'h34;
end 12'h1b6:    begin Red = 8'h61;    Green = 8'h70;    Blue = 8'h29;
end 12'h1b7:    begin Red = 8'h88;    Green = 8'ha0;    Blue = 8'h19;
end 12'h1b8:    begin Red = 8'h83;    Green = 8'h9a;    Blue = 8'h1b;
end 12'h1b9:    begin Red = 8'h3e;    Green = 8'h5f;    Blue = 8'h5f;
end 12'h1ba:    begin Red = 8'h5e;    Green = 8'h48;    Blue = 8'h34;
end 12'h1bb:    begin Red = 8'hd4;    Green = 8'hd2;    Blue = 8'hcf;
end 12'h1bc:    begin Red = 8'he3;    Green = 8'hd4;    Blue = 8'hc9;
end 12'h1bd:    begin Red = 8'h44;    Green = 8'h64;    Blue = 8'h46;
end 12'h1be:    begin Red = 8'hd7;    Green = 8'hda;    Blue = 8'hd1;
end 12'h1bf:    begin Red = 8'h49;    Green = 8'h59;    Blue = 8'h45;
end 12'h1c0:    begin Red = 8'hef;    Green = 8'he3;    Blue = 8'he3;
end 12'h1c1:    begin Red = 8'h4d;    Green = 8'h5e;    Blue = 8'h47;
end 12'h1c2:    begin Red = 8'h51;    Green = 8'h5c;    Blue = 8'h4c;
end 12'h1c3:    begin Red = 8'hcd;    Green = 8'hc7;    Blue = 8'hc3;
end 12'h1c4:    begin Red = 8'hcd;    Green = 8'hc6;    Blue = 8'h9d;
end 12'h1c5:    begin Red = 8'h02;    Green = 8'ha3;    Blue = 8'h3e;
end 12'h1c6:    begin Red = 8'h4e;    Green = 8'h59;    Blue = 8'h27;
end 12'h1c7:    begin Red = 8'h03;    Green = 8'h53;    Blue = 8'h79;
end 12'h1c8:    begin Red = 8'h02;    Green = 8'ha3;    Blue = 8'hfe;
end 12'h1c9:    begin Red = 8'h2d;    Green = 8'h36;    Blue = 8'h11;
end 12'h1ca:    begin Red = 8'h59;    Green = 8'h68;    Blue = 8'h21;
end 12'h1cb:    begin Red = 8'h55;    Green = 8'h63;    Blue = 8'h22;
end 12'h1cc:    begin Red = 8'h40;    Green = 8'h33;    Blue = 8'h36;
end 12'h1cd:    begin Red = 8'h47;    Green = 8'h43;    Blue = 8'h3d;
end 12'h1ce:    begin Red = 8'h60;    Green = 8'h6f;    Blue = 8'h30;
end 12'h1cf:    begin Red = 8'h09;    Green = 8'h2a;    Blue = 8'h99;
end 12'h1d0:    begin Red = 8'h09;    Green = 8'h2a;    Blue = 8'h80;
end 12'h1d1:    begin Red = 8'h0a;    Green = 8'h8c;    Blue = 8'h57;
end 12'h1d2:    begin Red = 8'h0b;    Green = 8'hdd;    Blue = 8'h40;
end 12'h1d3:    begin Red = 8'h7c;    Green = 8'h65;    Blue = 8'h3b;
end 12'h1d4:    begin Red = 8'h97;    Green = 8'h7e;    Blue = 8'h56;
end 12'h1d5:    begin Red = 8'h64;    Green = 8'h4a;    Blue = 8'h35;
end 12'h1d6:    begin Red = 8'h59;    Green = 8'h47;    Blue = 8'h2c;
end 12'h1d7:    begin Red = 8'hf4;    Green = 8'hd1;    Blue = 8'haa;
end 12'h1d8:    begin Red = 8'hf3;    Green = 8'hec;    Blue = 8'he6;
end 12'h1d9:    begin Red = 8'h7a;    Green = 8'ha0;    Blue = 8'h7b;
end 12'h1da:    begin Red = 8'h6a;    Green = 8'h91;    Blue = 8'h6d;
end 12'h1db:    begin Red = 8'h5f;    Green = 8'h8f;    Blue = 8'h5b;
end 12'h1dc:    begin Red = 8'h42;    Green = 8'h5f;    Blue = 8'h3a;
end 12'h1dd:    begin Red = 8'h55;    Green = 8'h62;    Blue = 8'h49;
end 12'h1de:    begin Red = 8'hfc;    Green = 8'he3;    Blue = 8'hea;
end 12'h1df:    begin Red = 8'hf3;    Green = 8'he9;    Blue = 8'hec;
end 12'h1e0:    begin Red = 8'hda;    Green = 8'hd4;    Blue = 8'hcc;
end 12'h1e1:    begin Red = 8'hcb;    Green = 8'hc5;    Blue = 8'hbd;
end 12'h1e2:    begin Red = 8'hc2;    Green = 8'hc6;    Blue = 8'hb6;
end 12'h1e3:    begin Red = 8'h4a;    Green = 8'h60;    Blue = 8'h4e;
end 12'h1e4:    begin Red = 8'hc2;    Green = 8'hcb;    Blue = 8'hb9;
end 12'h1e5:    begin Red = 8'h48;    Green = 8'h67;    Blue = 8'h3f;
end 12'h1e6:    begin Red = 8'h3a;    Green = 8'h5a;    Blue = 8'h3e;
end 12'h1e7:    begin Red = 8'hcb;    Green = 8'hc0;    Blue = 8'hbc;
end 12'h1e8:    begin Red = 8'h34;    Green = 8'h3b;    Blue = 8'h12;
end 12'h1e9:    begin Red = 8'h55;    Green = 8'h5b;    Blue = 8'h25;
end 12'h1ea:    begin Red = 8'h45;    Green = 8'h41;    Blue = 8'h2f;
end 12'h1eb:    begin Red = 8'h4b;    Green = 8'h4a;    Blue = 8'h26;
end 12'h1ec:    begin Red = 8'h08;    Green = 8'hba;    Blue = 8'h3f;
end 12'h1ed:    begin Red = 8'h7e;    Green = 8'h93;    Blue = 8'h12;
end 12'h1ee:    begin Red = 8'h94;    Green = 8'hae;    Blue = 8'h1e;
end 12'h1ef:    begin Red = 8'h0b;    Green = 8'h2c;    Blue = 8'h0a;
end 12'h1f0:    begin Red = 8'hb0;    Green = 8'h92;    Blue = 8'h69;
end 12'h1f1:    begin Red = 8'h44;    Green = 8'h59;    Blue = 8'h41;
end 12'h1f2:    begin Red = 8'h39;    Green = 8'h57;    Blue = 8'h4f;
end 12'h1f3:    begin Red = 8'hbd;    Green = 8'hb8;    Blue = 8'h96;
end 12'h1f4:    begin Red = 8'h6d;    Green = 8'h6e;    Blue = 8'h54;
end 12'h1f5:    begin Red = 8'h9d;    Green = 8'h9e;    Blue = 8'h88;
end 12'h1f6:    begin Red = 8'h98;    Green = 8'h9a;    Blue = 8'h81;
end 12'h1f7:    begin Red = 8'h03;    Green = 8'h23;    Blue = 8'hac;
end 12'h1f8:    begin Red = 8'h02;    Green = 8'hf3;    Blue = 8'h4e;
end 12'h1f9:    begin Red = 8'h02;    Green = 8'hf3;    Blue = 8'ha9;
end 12'h1fa:    begin Red = 8'h4d;    Green = 8'h4b;    Blue = 8'h36;
end 12'h1fb:    begin Red = 8'h4d;    Green = 8'h4b;    Blue = 8'h2b;
end 12'h1fc:    begin Red = 8'h46;    Green = 8'h49;    Blue = 8'h2d;
end 12'h1fd:    begin Red = 8'h61;    Green = 8'h76;    Blue = 8'h2b;
end 12'h1fe:    begin Red = 8'h6a;    Green = 8'h7a;    Blue = 8'h1c;
end 12'h1ff:    begin Red = 8'h3f;    Green = 8'h5e;    Blue = 8'h57;
end 12'h200:    begin Red = 8'h7b;    Green = 8'h95;    Blue = 8'h2e;
end 12'h201:    begin Red = 8'h7e;    Green = 8'ha9;    Blue = 8'h87;
end 12'h202:    begin Red = 8'hf1;    Green = 8'he4;    Blue = 8'hea;
end 12'h203:    begin Red = 8'hd1;    Green = 8'hda;    Blue = 8'hd1;
end 12'h204:    begin Red = 8'h4a;    Green = 8'h6a;    Blue = 8'h4d;
end 12'h205:    begin Red = 8'hc5;    Green = 8'hbf;    Blue = 8'hb8;
end 12'h206:    begin Red = 8'h76;    Green = 8'h71;    Blue = 8'h63;
end 12'h207:    begin Red = 8'h79;    Green = 8'h8a;    Blue = 8'h2e;
end 12'h208:    begin Red = 8'h9b;    Green = 8'h9a;    Blue = 8'h9b;
end 12'h209:    begin Red = 8'h02;    Green = 8'h62;    Blue = 8'hfe;
end 12'h20a:    begin Red = 8'h02;    Green = 8'h42;    Blue = 8'hdc;
end 12'h20b:    begin Red = 8'h55;    Green = 8'h5c;    Blue = 8'h32;
end 12'h20c:    begin Red = 8'h54;    Green = 8'h5b;    Blue = 8'h2a;
end 12'h20d:    begin Red = 8'h02;    Green = 8'he3;    Blue = 8'h53;
end 12'h20e:    begin Red = 8'h40;    Green = 8'h3c;    Blue = 8'h32;
end 12'h20f:    begin Red = 8'h71;    Green = 8'h74;    Blue = 8'h27;
end 12'h210:    begin Red = 8'h6d;    Green = 8'h87;    Blue = 8'h2a;
end 12'h211:    begin Red = 8'hba;    Green = 8'h9a;    Blue = 8'h7e;
end 12'h212:    begin Red = 8'hc4;    Green = 8'h93;    Blue = 8'h7d;
end 12'h213:    begin Red = 8'h70;    Green = 8'h50;    Blue = 8'h3d;
end 12'h214:    begin Red = 8'h6b;    Green = 8'h4b;    Blue = 8'h38;
end 12'h215:    begin Red = 8'h9e;    Green = 8'h7e;    Blue = 8'h66;
end 12'h216:    begin Red = 8'h97;    Green = 8'h77;    Blue = 8'h61;
end 12'h217:    begin Red = 8'hb1;    Green = 8'h8c;    Blue = 8'h77;
end 12'h218:    begin Red = 8'hb7;    Green = 8'h8c;    Blue = 8'h6c;
end 12'h219:    begin Red = 8'hcb;    Green = 8'ha3;    Blue = 8'h8b;
end 12'h21a:    begin Red = 8'h76;    Green = 8'h67;    Blue = 8'h3f;
end 12'h21b:    begin Red = 8'he9;    Green = 8'hd7;    Blue = 8'ha2;
end 12'h21c:    begin Red = 8'h98;    Green = 8'h75;    Blue = 8'h58;
end 12'h21d:    begin Red = 8'hfe;    Green = 8'he3;    Blue = 8'hc3;
end 12'h21e:    begin Red = 8'hff;    Green = 8'hec;    Blue = 8'hc0;
end 12'h21f:    begin Red = 8'h74;    Green = 8'h90;    Blue = 8'h36;
end 12'h220:    begin Red = 8'h7b;    Green = 8'h94;    Blue = 8'h33;
end 12'h221:    begin Red = 8'h87;    Green = 8'ha2;    Blue = 8'h8d;
end 12'h222:    begin Red = 8'hd9;    Green = 8'hce;    Blue = 8'hce;
end 12'h223:    begin Red = 8'h83;    Green = 8'h85;    Blue = 8'h67;
end 12'h224:    begin Red = 8'ha2;    Green = 8'h9e;    Blue = 8'h9e;
end 12'h225:    begin Red = 8'hb6;    Green = 8'hb2;    Blue = 8'hb3;
end 12'h226:    begin Red = 8'hb3;    Green = 8'haf;    Blue = 8'hae;
end 12'h227:    begin Red = 8'hab;    Green = 8'ha9;    Blue = 8'ha5;
end 12'h228:    begin Red = 8'h81;    Green = 8'h7b;    Blue = 8'h74;
end 12'h229:    begin Red = 8'h9a;    Green = 8'h94;    Blue = 8'ha9;
end 12'h22a:    begin Red = 8'h32;    Green = 8'h36;    Blue = 8'h20;
end 12'h22b:    begin Red = 8'h03;    Green = 8'h03;    Blue = 8'hbc;
end 12'h22c:    begin Red = 8'h3a;    Green = 8'h41;    Blue = 8'h1a;
end 12'h22d:    begin Red = 8'h29;    Green = 8'h31;    Blue = 8'h12;
end 12'h22e:    begin Red = 8'h61;    Green = 8'h62;    Blue = 8'h39;
end 12'h22f:    begin Red = 8'h5f;    Green = 8'h5e;    Blue = 8'h2b;
end 12'h230:    begin Red = 8'h62;    Green = 8'h5d;    Blue = 8'h36;
end 12'h231:    begin Red = 8'h38;    Green = 8'h57;    Blue = 8'h48;
end 12'h232:    begin Red = 8'hab;    Green = 8'h8e;    Blue = 8'h62;
end 12'h233:    begin Red = 8'h69;    Green = 8'h52;    Blue = 8'h43;
end 12'h234:    begin Red = 8'h75;    Green = 8'h55;    Blue = 8'h38;
end 12'h235:    begin Red = 8'h41;    Green = 8'h5e;    Blue = 8'h1e;
end 12'h236:    begin Red = 8'h3e;    Green = 8'h4f;    Blue = 8'h11;
end 12'h237:    begin Red = 8'hba;    Green = 8'h93;    Blue = 8'h7f;
end 12'h238:    begin Red = 8'hd4;    Green = 8'ha9;    Blue = 8'h90;
end 12'h239:    begin Red = 8'h7c;    Green = 8'h8d;    Blue = 8'h23;
end 12'h23a:    begin Red = 8'h72;    Green = 8'h94;    Blue = 8'h2b;
end 12'h23b:    begin Red = 8'h67;    Green = 8'h74;    Blue = 8'h59;
end 12'h23c:    begin Red = 8'h3f;    Green = 8'h66;    Blue = 8'h40;
end 12'h23d:    begin Red = 8'hc2;    Green = 8'hb8;    Blue = 8'hb2;
end 12'h23e:    begin Red = 8'hbc;    Green = 8'hb9;    Blue = 8'hb1;
end 12'h23f:    begin Red = 8'h66;    Green = 8'h7a;    Blue = 8'h51;
end 12'h240:    begin Red = 8'hb4;    Green = 8'hb4;    Blue = 8'h89;
end 12'h241:    begin Red = 8'h62;    Green = 8'h79;    Blue = 8'h19;
end 12'h242:    begin Red = 8'h72;    Green = 8'h75;    Blue = 8'h5a;
end 12'h243:    begin Red = 8'h04;    Green = 8'h75;    Blue = 8'h8e;
end 12'h244:    begin Red = 8'hb9;    Green = 8'haf;    Blue = 8'hb8;
end 12'h245:    begin Red = 8'h05;    Green = 8'h87;    Blue = 8'h1e;
end 12'h246:    begin Red = 8'h7a;    Green = 8'h96;    Blue = 8'h27;
end 12'h247:    begin Red = 8'h80;    Green = 8'h95;    Blue = 8'h3b;
end 12'h248:    begin Red = 8'h83;    Green = 8'h95;    Blue = 8'h36;
end 12'h249:    begin Red = 8'h99;    Green = 8'h99;    Blue = 8'h95;
end 12'h24a:    begin Red = 8'h67;    Green = 8'h76;    Blue = 8'h36;
end 12'h24b:    begin Red = 8'h4e;    Green = 8'h4d;    Blue = 8'h30;
end 12'h24c:    begin Red = 8'h47;    Green = 8'h3d;    Blue = 8'h35;
end 12'h24d:    begin Red = 8'h4e;    Green = 8'h45;    Blue = 8'h39;
end 12'h24e:    begin Red = 8'h53;    Green = 8'h4b;    Blue = 8'h40;
end 12'h24f:    begin Red = 8'h57;    Green = 8'h4d;    Blue = 8'h3b;
end 12'h250:    begin Red = 8'h6d;    Green = 8'h75;    Blue = 8'h31;
end 12'h251:    begin Red = 8'h66;    Green = 8'h59;    Blue = 8'h3e;
end 12'h252:    begin Red = 8'h9a;    Green = 8'h98;    Blue = 8'h1f;
end 12'h253:    begin Red = 8'h90;    Green = 8'h91;    Blue = 8'h27;
end 12'h254:    begin Red = 8'h96;    Green = 8'h91;    Blue = 8'h29;
end 12'h255:    begin Red = 8'h9b;    Green = 8'h8d;    Blue = 8'h1e;
end 12'h256:    begin Red = 8'h09;    Green = 8'h49;    Blue = 8'h5c;
end 12'h257:    begin Red = 8'hb8;    Green = 8'h97;    Blue = 8'h1b;
end 12'h258:    begin Red = 8'h78;    Green = 8'h5d;    Blue = 8'h43;
end 12'h259:    begin Red = 8'hbe;    Green = 8'h9f;    Blue = 8'h75;
end 12'h25a:    begin Red = 8'hc3;    Green = 8'ha5;    Blue = 8'h7c;
end 12'h25b:    begin Red = 8'hb2;    Green = 8'h9a;    Blue = 8'h73;
end 12'h25c:    begin Red = 8'h62;    Green = 8'h80;    Blue = 8'h22;
end 12'h25d:    begin Red = 8'h03;    Green = 8'hc4;    Blue = 8'h9e;
end 12'h25e:    begin Red = 8'h03;    Green = 8'he5;    Blue = 8'h2e;
end 12'h25f:    begin Red = 8'h72;    Green = 8'h80;    Blue = 8'h2c;
end 12'h260:    begin Red = 8'h79;    Green = 8'h7e;    Blue = 8'h33;
end 12'h261:    begin Red = 8'h33;    Green = 8'h4e;    Blue = 8'h13;
end 12'h262:    begin Red = 8'h03;    Green = 8'h84;    Blue = 8'hab;
end 12'h263:    begin Red = 8'h5e;    Green = 8'h6d;    Blue = 8'h24;
end 12'h264:    begin Red = 8'h54;    Green = 8'h6a;    Blue = 8'h18;
end 12'h265:    begin Red = 8'h02;    Green = 8'h53;    Blue = 8'hb0;
end 12'h266:    begin Red = 8'h04;    Green = 8'h15;    Blue = 8'h5b;
end 12'h267:    begin Red = 8'h02;    Green = 8'h44;    Blue = 8'h00;
end 12'h268:    begin Red = 8'h03;    Green = 8'h04;    Blue = 8'h42;
end 12'h269:    begin Red = 8'h4a;    Green = 8'h53;    Blue = 8'h14;
end 12'h26a:    begin Red = 8'h8d;    Green = 8'ha3;    Blue = 8'h31;
end 12'h26b:    begin Red = 8'h80;    Green = 8'ha8;    Blue = 8'h8f;
end 12'h26c:    begin Red = 8'h83;    Green = 8'ha2;    Blue = 8'h94;
end 12'h26d:    begin Red = 8'h82;    Green = 8'ha9;    Blue = 8'h7b;
end 12'h26e:    begin Red = 8'hce;    Green = 8'hd4;    Blue = 8'hd2;
end 12'h26f:    begin Red = 8'he1;    Green = 8'hd2;    Blue = 8'hd6;
end 12'h270:    begin Red = 8'heb;    Green = 8'hdb;    Blue = 8'he4;
end 12'h271:    begin Red = 8'hbf;    Green = 8'hc3;    Blue = 8'hbe;
end 12'h272:    begin Red = 8'h4b;    Green = 8'h5e;    Blue = 8'h41;
end 12'h273:    begin Red = 8'h66;    Green = 8'h6f;    Blue = 8'h64;
end 12'h274:    begin Red = 8'h39;    Green = 8'h4f;    Blue = 8'h5b;
end 12'h275:    begin Red = 8'hc3;    Green = 8'hbc;    Blue = 8'h93;
end 12'h276:    begin Red = 8'hb6;    Green = 8'hb4;    Blue = 8'h8f;
end 12'h277:    begin Red = 8'h63;    Green = 8'h70;    Blue = 8'h19;
end 12'h278:    begin Red = 8'h61;    Green = 8'h74;    Blue = 8'h1f;
end 12'h279:    begin Red = 8'h03;    Green = 8'hb4;    Blue = 8'h52;
end 12'h27a:    begin Red = 8'h03;    Green = 8'h04;    Blue = 8'h56;
end 12'h27b:    begin Red = 8'h5a;    Green = 8'h73;    Blue = 8'h2b;
end 12'h27c:    begin Red = 8'h53;    Green = 8'h72;    Blue = 8'h11;
end 12'h27d:    begin Red = 8'h03;    Green = 8'h94;    Blue = 8'he6;
end 12'h27e:    begin Red = 8'h86;    Green = 8'h9e;    Blue = 8'h30;
end 12'h27f:    begin Red = 8'h72;    Green = 8'h61;    Blue = 8'h60;
end 12'h280:    begin Red = 8'h61;    Green = 8'h5b;    Blue = 8'h5d;
end 12'h281:    begin Red = 8'h90;    Green = 8'h89;    Blue = 8'h8d;
end 12'h282:    begin Red = 8'h97;    Green = 8'h94;    Blue = 8'h8d;
end 12'h283:    begin Red = 8'h6b;    Green = 8'h75;    Blue = 8'h29;
end 12'h284:    begin Red = 8'h4a;    Green = 8'h44;    Blue = 8'h30;
end 12'h285:    begin Red = 8'h40;    Green = 8'h43;    Blue = 8'h2a;
end 12'h286:    begin Red = 8'h3e;    Green = 8'h3c;    Blue = 8'h37;
end 12'h287:    begin Red = 8'h37;    Green = 8'h36;    Blue = 8'h35;
end 12'h288:    begin Red = 8'h5d;    Green = 8'h69;    Blue = 8'h32;
end 12'h289:    begin Red = 8'h5f;    Green = 8'h4f;    Blue = 8'h3b;
end 12'h28a:    begin Red = 8'h9f;    Green = 8'h94;    Blue = 8'h20;
end 12'h28b:    begin Red = 8'h99;    Green = 8'h8f;    Blue = 8'h23;
end 12'h28c:    begin Red = 8'h93;    Green = 8'h87;    Blue = 8'h27;
end 12'h28d:    begin Red = 8'h8c;    Green = 8'h88;    Blue = 8'h24;
end 12'h28e:    begin Red = 8'h87;    Green = 8'h8b;    Blue = 8'h20;
end 12'h28f:    begin Red = 8'h9d;    Green = 8'h90;    Blue = 8'h13;
end 12'h290:    begin Red = 8'h21;    Green = 8'h46;    Blue = 8'h74;
end 12'h291:    begin Red = 8'h2c;    Green = 8'h4b;    Blue = 8'h6f;
end 12'h292:    begin Red = 8'hb4;    Green = 8'h98;    Blue = 8'h7d;
end 12'h293:    begin Red = 8'h50;    Green = 8'h74;    Blue = 8'h24;
end 12'h294:    begin Red = 8'h75;    Green = 8'h84;    Blue = 8'h3a;
end 12'h295:    begin Red = 8'h45;    Green = 8'h52;    Blue = 8'h15;
end 12'h296:    begin Red = 8'hff;    Green = 8'hfa;    Blue = 8'hcd;
end 12'h297:    begin Red = 8'h03;    Green = 8'h64;    Blue = 8'haf;
end 12'h298:    begin Red = 8'h48;    Green = 8'h55;    Blue = 8'h1a;
end 12'h299:    begin Red = 8'h59;    Green = 8'h6f;    Blue = 8'h1d;
end 12'h29a:    begin Red = 8'h04;    Green = 8'h76;    Blue = 8'h3a;
end 12'h29b:    begin Red = 8'h64;    Green = 8'h83;    Blue = 8'h16;
end 12'h29c:    begin Red = 8'h7d;    Green = 8'ha2;    Blue = 8'h81;
end 12'h29d:    begin Red = 8'h75;    Green = 8'h99;    Blue = 8'h70;
end 12'h29e:    begin Red = 8'hde;    Green = 8'he4;    Blue = 8'hde;
end 12'h29f:    begin Red = 8'h72;    Green = 8'h97;    Blue = 8'h69;
end 12'h2a0:    begin Red = 8'h44;    Green = 8'h6c;    Blue = 8'h43;
end 12'h2a1:    begin Red = 8'h3a;    Green = 8'h5d;    Blue = 8'h36;
end 12'h2a2:    begin Red = 8'hd8;    Green = 8'hc5;    Blue = 8'hc8;
end 12'h2a3:    begin Red = 8'h5c;    Green = 8'h6d;    Blue = 8'h51;
end 12'h2a4:    begin Red = 8'h4c;    Green = 8'h70;    Blue = 8'h43;
end 12'h2a5:    begin Red = 8'h63;    Green = 8'h79;    Blue = 8'h1f;
end 12'h2a6:    begin Red = 8'h42;    Green = 8'h4f;    Blue = 8'h1e;
end 12'h2a7:    begin Red = 8'h04;    Green = 8'h35;    Blue = 8'h1d;
end 12'h2a8:    begin Red = 8'h4c;    Green = 8'h55;    Blue = 8'h2f;
end 12'h2a9:    begin Red = 8'h05;    Green = 8'ha6;    Blue = 8'hde;
end 12'h2aa:    begin Red = 8'hc7;    Green = 8'hb6;    Blue = 8'hb7;
end 12'h2ab:    begin Red = 8'ha6;    Green = 8'hb0;    Blue = 8'ha8;
end 12'h2ac:    begin Red = 8'h5c;    Green = 8'h72;    Blue = 8'h24;
end 12'h2ad:    begin Red = 8'h6d;    Green = 8'h73;    Blue = 8'h52;
end 12'h2ae:    begin Red = 8'h5e;    Green = 8'h65;    Blue = 8'h54;
end 12'h2af:    begin Red = 8'h92;    Green = 8'h99;    Blue = 8'h91;
end 12'h2b0:    begin Red = 8'h49;    Green = 8'h46;    Blue = 8'h38;
end 12'h2b1:    begin Red = 8'h9c;    Green = 8'h93;    Blue = 8'h29;
end 12'h2b2:    begin Red = 8'h89;    Green = 8'h85;    Blue = 8'h1a;
end 12'h2b3:    begin Red = 8'h8b;    Green = 8'h7f;    Blue = 8'h25;
end 12'h2b4:    begin Red = 8'h7e;    Green = 8'h84;    Blue = 8'h24;
end 12'h2b5:    begin Red = 8'had;    Green = 8'haf;    Blue = 8'h1e;
end 12'h2b6:    begin Red = 8'ha2;    Green = 8'h91;    Blue = 8'h13;
end 12'h2b7:    begin Red = 8'h50;    Green = 8'h5f;    Blue = 8'h21;
end 12'h2b8:    begin Red = 8'h06;    Green = 8'h27;    Blue = 8'hde;
end 12'h2b9:    begin Red = 8'h70;    Green = 8'h98;    Blue = 8'h6e;
end 12'h2ba:    begin Red = 8'hc9;    Green = 8'hc8;    Blue = 8'hb6;
end 12'h2bb:    begin Red = 8'hc6;    Green = 8'hc5;    Blue = 8'hbb;
end 12'h2bc:    begin Red = 8'h66;    Green = 8'h80;    Blue = 8'h5d;
end 12'h2bd:    begin Red = 8'hb2;    Green = 8'hae;    Blue = 8'h85;
end 12'h2be:    begin Red = 8'h7b;    Green = 8'h7d;    Blue = 8'h60;
end 12'h2bf:    begin Red = 8'haa;    Green = 8'h74;    Blue = 8'h48;
end 12'h2c0:    begin Red = 8'ha0;    Green = 8'h6e;    Blue = 8'h42;
end 12'h2c1:    begin Red = 8'h81;    Green = 8'h89;    Blue = 8'h30;
end 12'h2c2:    begin Red = 8'h6e;    Green = 8'h68;    Blue = 8'h53;
end 12'h2c3:    begin Red = 8'h6c;    Green = 8'h75;    Blue = 8'h67;
end 12'h2c4:    begin Red = 8'h78;    Green = 8'h54;    Blue = 8'h33;
end 12'h2c5:    begin Red = 8'h8c;    Green = 8'h67;    Blue = 8'h44;
end 12'h2c6:    begin Red = 8'h5c;    Green = 8'h69;    Blue = 8'h2d;
end 12'h2c7:    begin Red = 8'h48;    Green = 8'h3e;    Blue = 8'h3e;
end 12'h2c8:    begin Red = 8'h68;    Green = 8'h71;    Blue = 8'h31;
end 12'h2c9:    begin Red = 8'h5d;    Green = 8'h55;    Blue = 8'h37;
end 12'h2ca:    begin Red = 8'h6e;    Green = 8'h57;    Blue = 8'h2d;
end 12'h2cb:    begin Red = 8'h6f;    Green = 8'h61;    Blue = 8'h2b;
end 12'h2cc:    begin Red = 8'h99;    Green = 8'h92;    Blue = 8'h1d;
end 12'h2cd:    begin Red = 8'h94;    Green = 8'h87;    Blue = 8'h1f;
end 12'h2ce:    begin Red = 8'h86;    Green = 8'h80;    Blue = 8'h2e;
end 12'h2cf:    begin Red = 8'hc2;    Green = 8'hb4;    Blue = 8'h2c;
end 12'h2d0:    begin Red = 8'h23;    Green = 8'h49;    Blue = 8'h65;
end 12'h2d1:    begin Red = 8'h24;    Green = 8'h4e;    Blue = 8'h5d;
end 12'h2d2:    begin Red = 8'hd9;    Green = 8'hb4;    Blue = 8'h8b;
end 12'h2d3:    begin Red = 8'hcb;    Green = 8'ha8;    Blue = 8'h86;
end 12'h2d4:    begin Red = 8'hfd;    Green = 8'hfc;    Blue = 8'hdd;
end 12'h2d5:    begin Red = 8'hfa;    Green = 8'hf1;    Blue = 8'hc9;
end 12'h2d6:    begin Red = 8'h78;    Green = 8'h8e;    Blue = 8'h15;
end 12'h2d7:    begin Red = 8'hff;    Green = 8'he1;    Blue = 8'hc8;
end 12'h2d8:    begin Red = 8'h7b;    Green = 8'ha1;    Blue = 8'h86;
end 12'h2d9:    begin Red = 8'h7f;    Green = 8'ha7;    Blue = 8'h81;
end 12'h2da:    begin Red = 8'he9;    Green = 8'hef;    Blue = 8'he5;
end 12'h2db:    begin Red = 8'hda;    Green = 8'he4;    Blue = 8'he7;
end 12'h2dc:    begin Red = 8'hda;    Green = 8'hd1;    Blue = 8'hd4;
end 12'h2dd:    begin Red = 8'hd5;    Green = 8'hdb;    Blue = 8'hd7;
end 12'h2de:    begin Red = 8'hd3;    Green = 8'hd9;    Blue = 8'hc9;
end 12'h2df:    begin Red = 8'hec;    Green = 8'he9;    Blue = 8'he4;
end 12'h2e0:    begin Red = 8'hd5;    Green = 8'hd5;    Blue = 8'hdb;
end 12'h2e1:    begin Red = 8'he5;    Green = 8'hd3;    Blue = 8'hd1;
end 12'h2e2:    begin Red = 8'hdb;    Green = 8'hd0;    Blue = 8'hdd;
end 12'h2e3:    begin Red = 8'hd0;    Green = 8'hc4;    Blue = 8'hb6;
end 12'h2e4:    begin Red = 8'h3e;    Green = 8'h55;    Blue = 8'h3c;
end 12'h2e5:    begin Red = 8'hb1;    Green = 8'hb6;    Blue = 8'haa;
end 12'h2e6:    begin Red = 8'h33;    Green = 8'h48;    Blue = 8'h30;
end 12'h2e7:    begin Red = 8'hbc;    Green = 8'hc4;    Blue = 8'hb8;
end 12'h2e8:    begin Red = 8'h2e;    Green = 8'h4a;    Blue = 8'h33;
end 12'h2e9:    begin Red = 8'h2e;    Green = 8'h47;    Blue = 8'h2d;
end 12'h2ea:    begin Red = 8'hbf;    Green = 8'hb3;    Blue = 8'had;
end 12'h2eb:    begin Red = 8'hc0;    Green = 8'hb6;    Blue = 8'h8e;
end 12'h2ec:    begin Red = 8'h72;    Green = 8'h82;    Blue = 8'h33;
end 12'h2ed:    begin Red = 8'hbc;    Green = 8'h7c;    Blue = 8'h5b;
end 12'h2ee:    begin Red = 8'hb5;    Green = 8'h7a;    Blue = 8'h47;
end 12'h2ef:    begin Red = 8'h5d;    Green = 8'h5a;    Blue = 8'h1d;
end 12'h2f0:    begin Red = 8'h60;    Green = 8'h5d;    Blue = 8'h24;
end 12'h2f1:    begin Red = 8'h58;    Green = 8'h64;    Blue = 8'h2b;
end 12'h2f2:    begin Red = 8'h69;    Green = 8'h61;    Blue = 8'h66;
end 12'h2f3:    begin Red = 8'h65;    Green = 8'h69;    Blue = 8'h69;
end 12'h2f4:    begin Red = 8'h8c;    Green = 8'h6b;    Blue = 8'h39;
end 12'h2f5:    begin Red = 8'h88;    Green = 8'h61;    Blue = 8'h39;
end 12'h2f6:    begin Red = 8'ha2;    Green = 8'hc1;    Blue = 8'h13;
end 12'h2f7:    begin Red = 8'h62;    Green = 8'h7d;    Blue = 8'h32;
end 12'h2f8:    begin Red = 8'h83;    Green = 8'h9b;    Blue = 8'h14;
end 12'h2f9:    begin Red = 8'h5f;    Green = 8'h6a;    Blue = 8'h37;
end 12'h2fa:    begin Red = 8'h08;    Green = 8'h59;    Blue = 8'hff;
end 12'h2fb:    begin Red = 8'h78;    Green = 8'h76;    Blue = 8'h24;
end 12'h2fc:    begin Red = 8'h71;    Green = 8'h5d;    Blue = 8'h32;
end 12'h2fd:    begin Red = 8'h61;    Green = 8'h5f;    Blue = 8'h30;
end 12'h2fe:    begin Red = 8'h84;    Green = 8'h89;    Blue = 8'h2b;
end 12'h2ff:    begin Red = 8'hb8;    Green = 8'had;    Blue = 8'h2b;
end 12'h300:    begin Red = 8'hb8;    Green = 8'ha7;    Blue = 8'h2b;
end 12'h301:    begin Red = 8'hb5;    Green = 8'haa;    Blue = 8'h35;
end 12'h302:    begin Red = 8'ha0;    Green = 8'h83;    Blue = 8'h72;
end 12'h303:    begin Red = 8'h94;    Green = 8'h89;    Blue = 8'h6a;
end 12'h304:    begin Red = 8'h1c;    Green = 8'h4a;    Blue = 8'h58;
end 12'h305:    begin Red = 8'h78;    Green = 8'h63;    Blue = 8'h49;
end 12'h306:    begin Red = 8'h6d;    Green = 8'h5c;    Blue = 8'h37;
end 12'h307:    begin Red = 8'h02;    Green = 8'h93;    Blue = 8'h39;
end 12'h308:    begin Red = 8'h03;    Green = 8'h13;    Blue = 8'hb2;
end 12'h309:    begin Red = 8'h40;    Green = 8'h4e;    Blue = 8'h17;
end 12'h30a:    begin Red = 8'h08;    Green = 8'h4a;    Blue = 8'h0f;
end 12'h30b:    begin Red = 8'h88;    Green = 8'h9b;    Blue = 8'h93;
end 12'h30c:    begin Red = 8'h74;    Green = 8'haa;    Blue = 8'h82;
end 12'h30d:    begin Red = 8'ha1;    Green = 8'h85;    Blue = 8'h64;
end 12'h30e:    begin Red = 8'h9d;    Green = 8'h8a;    Blue = 8'h6a;
end 12'h30f:    begin Red = 8'h92;    Green = 8'h90;    Blue = 8'h8b;
end 12'h310:    begin Red = 8'he7;    Green = 8'hdb;    Blue = 8'hde;
end 12'h311:    begin Red = 8'hbe;    Green = 8'hc5;    Blue = 8'hb0;
end 12'h312:    begin Red = 8'h96;    Green = 8'h8f;    Blue = 8'h90;
end 12'h313:    begin Red = 8'h8b;    Green = 8'h90;    Blue = 8'h85;
end 12'h314:    begin Red = 8'ha8;    Green = 8'h91;    Blue = 8'h8b;
end 12'h315:    begin Red = 8'hd9;    Green = 8'hcc;    Blue = 8'hc1;
end 12'h316:    begin Red = 8'hc0;    Green = 8'hbc;    Blue = 8'hb9;
end 12'h317:    begin Red = 8'hb3;    Green = 8'had;    Blue = 8'ha6;
end 12'h318:    begin Red = 8'hb9;    Green = 8'had;    Blue = 8'haa;
end 12'h319:    begin Red = 8'h70;    Green = 8'h7b;    Blue = 8'h53;
end 12'h31a:    begin Red = 8'h62;    Green = 8'h76;    Blue = 8'h32;
end 12'h31b:    begin Red = 8'h03;    Green = 8'h13;    Blue = 8'h9e;
end 12'h31c:    begin Red = 8'h03;    Green = 8'h43;    Blue = 8'hce;
end 12'h31d:    begin Red = 8'h4d;    Green = 8'h5d;    Blue = 8'h16;
end 12'h31e:    begin Red = 8'h02;    Green = 8'h93;    Blue = 8'h4d;
end 12'h31f:    begin Red = 8'h57;    Green = 8'h6b;    Blue = 8'h26;
end 12'h320:    begin Red = 8'h02;    Green = 8'he3;    Blue = 8'h4c;
end 12'h321:    begin Red = 8'h41;    Green = 8'h2d;    Blue = 8'h34;
end 12'h322:    begin Red = 8'h07;    Green = 8'hb9;    Blue = 8'hfe;
end 12'h323:    begin Red = 8'h73;    Green = 8'h52;    Blue = 8'h2b;
end 12'h324:    begin Red = 8'h88;    Green = 8'ha1;    Blue = 8'h13;
end 12'h325:    begin Red = 8'h7e;    Green = 8'h94;    Blue = 8'h1d;
end 12'h326:    begin Red = 8'h09;    Green = 8'h8a;    Blue = 8'h24;
end 12'h327:    begin Red = 8'h99;    Green = 8'h83;    Blue = 8'h33;
end 12'h328:    begin Red = 8'h8c;    Green = 8'h84;    Blue = 8'h2a;
end 12'h329:    begin Red = 8'h9f;    Green = 8'h88;    Blue = 8'h73;
end 12'h32a:    begin Red = 8'h20;    Green = 8'h4f;    Blue = 8'h51;
end 12'h32b:    begin Red = 8'h7a;    Green = 8'h69;    Blue = 8'h4d;
end 12'h32c:    begin Red = 8'hcd;    Green = 8'had;    Blue = 8'h84;
end 12'h32d:    begin Red = 8'h03;    Green = 8'h33;    Blue = 8'h9f;
end 12'h32e:    begin Red = 8'h03;    Green = 8'h23;    Blue = 8'hba;
end 12'h32f:    begin Red = 8'h54;    Green = 8'h63;    Blue = 8'h1a;
end 12'h330:    begin Red = 8'h40;    Green = 8'h41;    Blue = 8'h32;
end 12'h331:    begin Red = 8'h9c;    Green = 8'hb9;    Blue = 8'h17;
end 12'h332:    begin Red = 8'h09;    Green = 8'hab;    Blue = 8'h80;
end 12'h333:    begin Red = 8'h9b;    Green = 8'h87;    Blue = 8'h64;
end 12'h334:    begin Red = 8'h80;    Green = 8'h89;    Blue = 8'h7f;
end 12'h335:    begin Red = 8'h95;    Green = 8'h88;    Blue = 8'h8d;
end 12'h336:    begin Red = 8'h85;    Green = 8'h8a;    Blue = 8'h80;
end 12'h337:    begin Red = 8'h89;    Green = 8'h81;    Blue = 8'h85;
end 12'h338:    begin Red = 8'h89;    Green = 8'h82;    Blue = 8'h8c;
end 12'h339:    begin Red = 8'h86;    Green = 8'h88;    Blue = 8'h86;
end 12'h33a:    begin Red = 8'h71;    Green = 8'h7d;    Blue = 8'h73;
end 12'h33b:    begin Red = 8'h7a;    Green = 8'h7b;    Blue = 8'h73;
end 12'h33c:    begin Red = 8'h51;    Green = 8'h5d;    Blue = 8'h52;
end 12'h33d:    begin Red = 8'h43;    Green = 8'h5e;    Blue = 8'h47;
end 12'h33e:    begin Red = 8'ha7;    Green = 8'ha8;    Blue = 8'h86;
end 12'h33f:    begin Red = 8'h30;    Green = 8'h35;    Blue = 8'h1b;
end 12'h340:    begin Red = 8'h02;    Green = 8'h83;    Blue = 8'h6f;
end 12'h341:    begin Red = 8'h3d;    Green = 8'h3a;    Blue = 8'h13;
end 12'h342:    begin Red = 8'h5a;    Green = 8'h6e;    Blue = 8'h34;
end 12'h343:    begin Red = 8'h9b;    Green = 8'hb3;    Blue = 8'h1d;
end 12'h344:    begin Red = 8'h95;    Green = 8'hb2;    Blue = 8'h18;
end 12'h345:    begin Red = 8'h08;    Green = 8'haa;    Blue = 8'h6a;
end 12'h346:    begin Red = 8'h93;    Green = 8'haf;    Blue = 8'h10;
end 12'h347:    begin Red = 8'h08;    Green = 8'h9a;    Blue = 8'h4e;
end 12'h348:    begin Red = 8'h09;    Green = 8'heb;    Blue = 8'hf5;
end 12'h349:    begin Red = 8'h3c;    Green = 8'h60;    Blue = 8'h78;
end 12'h34a:    begin Red = 8'h23;    Green = 8'h49;    Blue = 8'h56;
end 12'h34b:    begin Red = 8'h17;    Green = 8'h46;    Blue = 8'h5a;
end 12'h34c:    begin Red = 8'h0c;    Green = 8'h44;    Blue = 8'h5f;
end 12'h34d:    begin Red = 8'h87;    Green = 8'h8a;    Blue = 8'h15;
end 12'h34e:    begin Red = 8'h97;    Green = 8'h88;    Blue = 8'h75;
end 12'h34f:    begin Red = 8'h17;    Green = 8'h41;    Blue = 8'h52;
end 12'h350:    begin Red = 8'h5d;    Green = 8'h40;    Blue = 8'h31;
end 12'h351:    begin Red = 8'h5b;    Green = 8'h41;    Blue = 8'h2c;
end 12'h352:    begin Red = 8'h37;    Green = 8'h5c;    Blue = 8'h11;
end 12'h353:    begin Red = 8'h51;    Green = 8'h73;    Blue = 8'h17;
end 12'h354:    begin Red = 8'h03;    Green = 8'h13;    Blue = 8'h8f;
end 12'h355:    begin Red = 8'h46;    Green = 8'h3b;    Blue = 8'h2e;
end 12'h356:    begin Red = 8'h3a;    Green = 8'h2f;    Blue = 8'h2f;
end 12'h357:    begin Red = 8'h53;    Green = 8'h6a;    Blue = 8'h2d;
end 12'h358:    begin Red = 8'h08;    Green = 8'h99;    Blue = 8'hfb;
end 12'h359:    begin Red = 8'h07;    Green = 8'h59;    Blue = 8'h9a;
end 12'h35a:    begin Red = 8'h08;    Green = 8'heb;    Blue = 8'h7a;
end 12'h35b:    begin Red = 8'h08;    Green = 8'h0b;    Blue = 8'h03;
end 12'h35c:    begin Red = 8'h71;    Green = 8'h9a;    Blue = 8'h7a;
end 12'h35d:    begin Red = 8'h67;    Green = 8'ha7;    Blue = 8'h75;
end 12'h35e:    begin Red = 8'h81;    Green = 8'h7c;    Blue = 8'h8f;
end 12'h35f:    begin Red = 8'h6d;    Green = 8'h9d;    Blue = 8'h75;
end 12'h360:    begin Red = 8'h6f;    Green = 8'h84;    Blue = 8'h7f;
end 12'h361:    begin Red = 8'h6c;    Green = 8'h95;    Blue = 8'h77;
end 12'h362:    begin Red = 8'h8d;    Green = 8'h9f;    Blue = 8'h81;
end 12'h363:    begin Red = 8'h94;    Green = 8'h84;    Blue = 8'h87;
end 12'h364:    begin Red = 8'h58;    Green = 8'h73;    Blue = 8'h4b;
end 12'h365:    begin Red = 8'h8b;    Green = 8'h88;    Blue = 8'h81;
end 12'h366:    begin Red = 8'h81;    Green = 8'h81;    Blue = 8'h80;
end 12'h367:    begin Red = 8'h52;    Green = 8'h70;    Blue = 8'h4e;
end 12'h368:    begin Red = 8'he8;    Green = 8'hd6;    Blue = 8'hdb;
end 12'h369:    begin Red = 8'h81;    Green = 8'h7c;    Blue = 8'h7a;
end 12'h36a:    begin Red = 8'h85;    Green = 8'h7c;    Blue = 8'h87;
end 12'h36b:    begin Red = 8'hd5;    Green = 8'hc9;    Blue = 8'hcf;
end 12'h36c:    begin Red = 8'hcb;    Green = 8'hbb;    Blue = 8'hb6;
end 12'h36d:    begin Red = 8'h51;    Green = 8'h7c;    Blue = 8'h5f;
end 12'h36e:    begin Red = 8'h4c;    Green = 8'h70;    Blue = 8'h5d;
end 12'h36f:    begin Red = 8'h11;    Green = 8'h3f;    Blue = 8'h57;
end 12'h370:    begin Red = 8'had;    Green = 8'hb6;    Blue = 8'h93;
end 12'h371:    begin Red = 8'h03;    Green = 8'h34;    Blue = 8'h47;
end 12'h372:    begin Red = 8'h04;    Green = 8'h05;    Blue = 8'h3d;
end 12'h373:    begin Red = 8'h70;    Green = 8'h82;    Blue = 8'h16;
end 12'h374:    begin Red = 8'h02;    Green = 8'h73;    Blue = 8'h0c;
end 12'h375:    begin Red = 8'h50;    Green = 8'h6a;    Blue = 8'h1d;
end 12'h376:    begin Red = 8'h4f;    Green = 8'h62;    Blue = 8'h1b;
end 12'h377:    begin Red = 8'h42;    Green = 8'h41;    Blue = 8'h38;
end 12'h378:    begin Red = 8'h49;    Green = 8'h69;    Blue = 8'h1a;
end 12'h379:    begin Red = 8'h46;    Green = 8'h61;    Blue = 8'h24;
end 12'h37a:    begin Red = 8'h06;    Green = 8'he9;    Blue = 8'h5a;
end 12'h37b:    begin Red = 8'h08;    Green = 8'h5b;    Blue = 8'h4c;
end 12'h37c:    begin Red = 8'h08;    Green = 8'h5b;    Blue = 8'h64;
end 12'h37d:    begin Red = 8'h27;    Green = 8'h24;    Blue = 8'h1c;
end 12'h37e:    begin Red = 8'hf9;    Green = 8'hd8;    Blue = 8'h9e;
end 12'h37f:    begin Red = 8'he7;    Green = 8'hbe;    Blue = 8'h9c;
end 12'h380:    begin Red = 8'ha6;    Green = 8'h83;    Blue = 8'h65;
end 12'h381:    begin Red = 8'hbb;    Green = 8'haa;    Blue = 8'h7d;
end 12'h382:    begin Red = 8'hfa;    Green = 8'hdd;    Blue = 8'hbb;
end 12'h383:    begin Red = 8'h73;    Green = 8'h57;    Blue = 8'h41;
end 12'h384:    begin Red = 8'h03;    Green = 8'h84;    Blue = 8'h9f;
end 12'h385:    begin Red = 8'h03;    Green = 8'h03;    Blue = 8'h6b;
end 12'h386:    begin Red = 8'hde;    Green = 8'hc0;    Blue = 8'h96;
end 12'h387:    begin Red = 8'hd8;    Green = 8'hb9;    Blue = 8'h98;
end 12'h388:    begin Red = 8'hdc;    Green = 8'hb9;    Blue = 8'h89;
end 12'h389:    begin Red = 8'he7;    Green = 8'hc8;    Blue = 8'h99;
end 12'h38a:    begin Red = 8'hba;    Green = 8'ha4;    Blue = 8'h7d;
end 12'h38b:    begin Red = 8'h82;    Green = 8'h84;    Blue = 8'h7a;
end 12'h38c:    begin Red = 8'h87;    Green = 8'h7b;    Blue = 8'h7c;
end 12'h38d:    begin Red = 8'h90;    Green = 8'h85;    Blue = 8'h82;
end 12'h38e:    begin Red = 8'h87;    Green = 8'h7c;    Blue = 8'h81;
end 12'h38f:    begin Red = 8'h77;    Green = 8'h70;    Blue = 8'h6f;
end 12'h390:    begin Red = 8'h9d;    Green = 8'h7c;    Blue = 8'h51;
end 12'h391:    begin Red = 8'hd9;    Green = 8'hae;    Blue = 8'h7e;
end 12'h392:    begin Red = 8'hd4;    Green = 8'h9d;    Blue = 8'h69;
end 12'h393:    begin Red = 8'hcd;    Green = 8'h9a;    Blue = 8'h6d;
end 12'h394:    begin Red = 8'hc9;    Green = 8'h9f;    Blue = 8'h69;
end 12'h395:    begin Red = 8'hce;    Green = 8'h98;    Blue = 8'h67;
end 12'h396:    begin Red = 8'h86;    Green = 8'h4f;    Blue = 8'h29;
end 12'h397:    begin Red = 8'h89;    Green = 8'h64;    Blue = 8'h33;
end 12'h398:    begin Red = 8'h71;    Green = 8'h6c;    Blue = 8'h66;
end 12'h399:    begin Red = 8'hce;    Green = 8'ha0;    Blue = 8'h6d;
end 12'h39a:    begin Red = 8'h65;    Green = 8'h5e;    Blue = 8'h2b;
end 12'h39b:    begin Red = 8'h53;    Green = 8'h4b;    Blue = 8'h30;
end 12'h39c:    begin Red = 8'h8e;    Green = 8'ha3;    Blue = 8'h15;
end 12'h39d:    begin Red = 8'h08;    Green = 8'h6a;    Blue = 8'h0e;
end 12'h39e:    begin Red = 8'h08;    Green = 8'h6a;    Blue = 8'h1b;
end 12'h39f:    begin Red = 8'h08;    Green = 8'hca;    Blue = 8'h8a;
end 12'h3a0:    begin Red = 8'h9c;    Green = 8'hb6;    Blue = 8'h24;
end 12'h3a1:    begin Red = 8'h00;    Green = 8'h0b;    Blue = 8'hfe;
end 12'h3a2:    begin Red = 8'h2f;    Green = 8'h35;    Blue = 8'h16;
end 12'h3a3:    begin Red = 8'h02;    Green = 8'hc3;    Blue = 8'h3e;
end 12'h3a4:    begin Red = 8'h03;    Green = 8'h84;    Blue = 8'hb7;
end 12'h3a5:    begin Red = 8'h03;    Green = 8'h33;    Blue = 8'hfa;
end 12'h3a6:    begin Red = 8'h02;    Green = 8'hb3;    Blue = 8'h86;
end 12'h3a7:    begin Red = 8'h9d;    Green = 8'h7f;    Blue = 8'h5d;
end 12'h3a8:    begin Red = 8'hda;    Green = 8'hbe;    Blue = 8'h8a;
end 12'h3a9:    begin Red = 8'hd4;    Green = 8'haf;    Blue = 8'h84;
end 12'h3aa:    begin Red = 8'hbf;    Green = 8'h98;    Blue = 8'h82;
end 12'h3ab:    begin Red = 8'h2a;    Green = 8'h38;    Blue = 8'h17;
end 12'h3ac:    begin Red = 8'h27;    Green = 8'h2c;    Blue = 8'h17;
end 12'h3ad:    begin Red = 8'h02;    Green = 8'h73;    Blue = 8'h2b;
end 12'h3ae:    begin Red = 8'h35;    Green = 8'h40;    Blue = 8'h12;
end 12'h3af:    begin Red = 8'h6c;    Green = 8'h81;    Blue = 8'h2d;
end 12'h3b0:    begin Red = 8'h66;    Green = 8'h57;    Blue = 8'h39;
end 12'h3b1:    begin Red = 8'h59;    Green = 8'h54;    Blue = 8'h27;
end 12'h3b2:    begin Red = 8'h5d;    Green = 8'h5a;    Blue = 8'h33;
end 12'h3b3:    begin Red = 8'hd7;    Green = 8'hbb;    Blue = 8'h9e;
end 12'h3b4:    begin Red = 8'h7a;    Green = 8'h84;    Blue = 8'h7b;
end 12'h3b5:    begin Red = 8'h58;    Green = 8'h79;    Blue = 8'h56;
end 12'h3b6:    begin Red = 8'h4e;    Green = 8'h59;    Blue = 8'h42;
end 12'h3b7:    begin Red = 8'h3e;    Green = 8'h58;    Blue = 8'h34;
end 12'h3b8:    begin Red = 8'h97;    Green = 8'h89;    Blue = 8'h88;
end 12'h3b9:    begin Red = 8'h54;    Green = 8'h78;    Blue = 8'h64;
end 12'h3ba:    begin Red = 8'h7c;    Green = 8'h58;    Blue = 8'h22;
end 12'h3bb:    begin Red = 8'h88;    Green = 8'h56;    Blue = 8'h2b;
end 12'h3bc:    begin Red = 8'he7;    Green = 8'hab;    Blue = 8'h77;
end 12'h3bd:    begin Red = 8'hdb;    Green = 8'hac;    Blue = 8'h6f;
end 12'h3be:    begin Red = 8'he3;    Green = 8'ha5;    Blue = 8'h6d;
end 12'h3bf:    begin Red = 8'he1;    Green = 8'hae;    Blue = 8'h6a;
end 12'h3c0:    begin Red = 8'hf1;    Green = 8'hb3;    Blue = 8'h7d;
end 12'h3c1:    begin Red = 8'h82;    Green = 8'h92;    Blue = 8'h2e;
end 12'h3c2:    begin Red = 8'h2e;    Green = 8'h31;    Blue = 8'h10;
end 12'h3c3:    begin Red = 8'h02;    Green = 8'hf3;    Blue = 8'h9f;
end 12'h3c4:    begin Red = 8'h03;    Green = 8'h44;    Blue = 8'h0c;
end 12'h3c5:    begin Red = 8'h02;    Green = 8'hb3;    Blue = 8'h6e;
end 12'h3c6:    begin Red = 8'h03;    Green = 8'h63;    Blue = 8'hea;
end 12'h3c7:    begin Red = 8'h58;    Green = 8'h57;    Blue = 8'h32;
end 12'h3c8:    begin Red = 8'h60;    Green = 8'h5b;    Blue = 8'h3d;
end 12'h3c9:    begin Red = 8'h63;    Green = 8'h56;    Blue = 8'h2d;
end 12'h3ca:    begin Red = 8'h49;    Green = 8'h4e;    Blue = 8'h31;
end 12'h3cb:    begin Red = 8'h32;    Green = 8'h48;    Blue = 8'h1c;
end 12'h3cc:    begin Red = 8'hd9;    Green = 8'h9d;    Blue = 8'h6d;
end 12'h3cd:    begin Red = 8'h68;    Green = 8'h5e;    Blue = 8'h32;
end 12'h3ce:    begin Red = 8'h86;    Green = 8'h94;    Blue = 8'h19;
end 12'h3cf:    begin Red = 8'h69;    Green = 8'h7b;    Blue = 8'h22;
end 12'h3d0:    begin Red = 8'h57;    Green = 8'h62;    Blue = 8'h31;
end 12'h3d1:    begin Red = 8'h98;    Green = 8'hb1;    Blue = 8'h27;
end 12'h3d2:    begin Red = 8'h1b;    Green = 8'h21;    Blue = 8'h14;
end 12'h3d3:    begin Red = 8'h47;    Green = 8'h60;    Blue = 8'h1f;
end 12'h3d4:    begin Red = 8'h42;    Green = 8'h4a;    Blue = 8'h11;
end 12'h3d5:    begin Red = 8'ha5;    Green = 8'h7f;    Blue = 8'h60;
end 12'h3d6:    begin Red = 8'hc0;    Green = 8'ha6;    Blue = 8'h74;
end 12'h3d7:    begin Red = 8'ha3;    Green = 8'h92;    Blue = 8'h6f;
end 12'h3d8:    begin Red = 8'h03;    Green = 8'h13;    Blue = 8'h7e;
end 12'h3d9:    begin Red = 8'h39;    Green = 8'h3c;    Blue = 8'h1b;
end 12'h3da:    begin Red = 8'hc7;    Green = 8'h9e;    Blue = 8'h75;
end 12'h3db:    begin Red = 8'hda;    Green = 8'hb7;    Blue = 8'h93;
end 12'h3dc:    begin Red = 8'hd2;    Green = 8'hb7;    Blue = 8'h95;
end 12'h3dd:    begin Red = 8'h80;    Green = 8'h79;    Blue = 8'h80;
end 12'h3de:    begin Red = 8'h7a;    Green = 8'h7f;    Blue = 8'h78;
end 12'h3df:    begin Red = 8'h4a;    Green = 8'h54;    Blue = 8'h43;
end 12'h3e0:    begin Red = 8'h44;    Green = 8'h54;    Blue = 8'h40;
end 12'h3e1:    begin Red = 8'h7d;    Green = 8'h57;    Blue = 8'h2c;
end 12'h3e2:    begin Red = 8'h7e;    Green = 8'h5d;    Blue = 8'h2b;
end 12'h3e3:    begin Red = 8'hd2;    Green = 8'h9f;    Blue = 8'h63;
end 12'h3e4:    begin Red = 8'hc4;    Green = 8'ha2;    Blue = 8'h65;
end 12'h3e5:    begin Red = 8'h02;    Green = 8'hf3;    Blue = 8'hfc;
end 12'h3e6:    begin Red = 8'h03;    Green = 8'h33;    Blue = 8'hbd;
end 12'h3e7:    begin Red = 8'h67;    Green = 8'h78;    Blue = 8'h3b;
end 12'h3e8:    begin Red = 8'h40;    Green = 8'h50;    Blue = 8'h26;
end 12'h3e9:    begin Red = 8'hd3;    Green = 8'h99;    Blue = 8'h72;
end 12'h3ea:    begin Red = 8'hcf;    Green = 8'h9e;    Blue = 8'h68;
end 12'h3eb:    begin Red = 8'h45;    Green = 8'h3e;    Blue = 8'h28;
end 12'h3ec:    begin Red = 8'h4c;    Green = 8'h3a;    Blue = 8'h26;
end 12'h3ed:    begin Red = 8'h09;    Green = 8'heb;    Blue = 8'hae;
end 12'h3ee:    begin Red = 8'h9f;    Green = 8'hbd;    Blue = 8'h1d;
end 12'h3ef:    begin Red = 8'h3d;    Green = 8'h37;    Blue = 8'h1a;
end 12'h3f0:    begin Red = 8'h2d;    Green = 8'h3b;    Blue = 8'h10;
end 12'h3f1:    begin Red = 8'ha7;    Green = 8'h87;    Blue = 8'h6d;
end 12'h3f2:    begin Red = 8'h93;    Green = 8'h90;    Blue = 8'h1d;
end 12'h3f3:    begin Red = 8'h6b;    Green = 8'h56;    Blue = 8'h3a;
end 12'h3f4:    begin Red = 8'h91;    Green = 8'h7c;    Blue = 8'h59;
end 12'h3f5:    begin Red = 8'h77;    Green = 8'haa;    Blue = 8'h7c;
end 12'h3f6:    begin Red = 8'h87;    Green = 8'h81;    Blue = 8'h7b;
end 12'h3f7:    begin Red = 8'h5e;    Green = 8'h7c;    Blue = 8'h69;
end 12'h3f8:    begin Red = 8'h8d;    Green = 8'h8a;    Blue = 8'h1f;
end 12'h3f9:    begin Red = 8'h6a;    Green = 8'h9d;    Blue = 8'h58;
end 12'h3fa:    begin Red = 8'h6a;    Green = 8'h9a;    Blue = 8'h5e;
end 12'h3fb:    begin Red = 8'h6a;    Green = 8'h80;    Blue = 8'h26;
end 12'h3fc:    begin Red = 8'h43;    Green = 8'h31;    Blue = 8'h27;
end 12'h3fd:    begin Red = 8'h35;    Green = 8'h26;    Blue = 8'h2a;
end 12'h3fe:    begin Red = 8'h46;    Green = 8'h42;    Blue = 8'h23;
end 12'h3ff:    begin Red = 8'ha5;    Green = 8'hc2;    Blue = 8'h1f;
end 12'h400:    begin Red = 8'h40;    Green = 8'h27;    Blue = 8'h29;
end 12'h401:    begin Red = 8'h09;    Green = 8'h4b;    Blue = 8'h3c;
end 12'h402:    begin Red = 8'h43;    Green = 8'h37;    Blue = 8'h1b;
end 12'h403:    begin Red = 8'h79;    Green = 8'h6a;    Blue = 8'h38;
end 12'h404:    begin Red = 8'h02;    Green = 8'h93;    Blue = 8'h2e;
end 12'h405:    begin Red = 8'h5b;    Green = 8'h6f;    Blue = 8'h14;
end 12'h406:    begin Red = 8'h45;    Green = 8'h72;    Blue = 8'h18;
end 12'h407:    begin Red = 8'h08;    Green = 8'h98;    Blue = 8'h9f;
end 12'h408:    begin Red = 8'h94;    Green = 8'h8d;    Blue = 8'h18;
end 12'h409:    begin Red = 8'hac;    Green = 8'hd4;    Blue = 8'h13;
end 12'h40a:    begin Red = 8'h9f;    Green = 8'hc9;    Blue = 8'h13;
end 12'h40b:    begin Red = 8'h09;    Green = 8'h9c;    Blue = 8'h80;
end 12'h40c:    begin Red = 8'h73;    Green = 8'h87;    Blue = 8'h20;
end 12'h40d:    begin Red = 8'h71;    Green = 8'h89;    Blue = 8'h25;
end 12'h40e:    begin Red = 8'h87;    Green = 8'ha3;    Blue = 8'h20;
end 12'h40f:    begin Red = 8'h08;    Green = 8'h9a;    Blue = 8'hbb;
end 12'h410:    begin Red = 8'h57;    Green = 8'h54;    Blue = 8'h2d;
end 12'h411:    begin Red = 8'hc5;    Green = 8'hbb;    Blue = 8'h2c;
end 12'h412:    begin Red = 8'h82;    Green = 8'h7f;    Blue = 8'h18;
end 12'h413:    begin Red = 8'h88;    Green = 8'h83;    Blue = 8'h15;
end 12'h414:    begin Red = 8'ha1;    Green = 8'h8d;    Blue = 8'h64;
end 12'h415:    begin Red = 8'hb9;    Green = 8'hb5;    Blue = 8'hc6;
end 12'h416:    begin Red = 8'hae;    Green = 8'ha4;    Blue = 8'had;
end 12'h417:    begin Red = 8'h90;    Green = 8'ha5;    Blue = 8'h86;
end 12'h418:    begin Red = 8'h69;    Green = 8'h72;    Blue = 8'h1c;
end 12'h419:    begin Red = 8'h69;    Green = 8'h78;    Blue = 8'h16;
end 12'h41a:    begin Red = 8'h88;    Green = 8'h98;    Blue = 8'h29;
end 12'h41b:    begin Red = 8'h66;    Green = 8'h71;    Blue = 8'h25;
end 12'h41c:    begin Red = 8'h7a;    Green = 8'h95;    Blue = 8'h22;
end 12'h41d:    begin Red = 8'h75;    Green = 8'h95;    Blue = 8'h26;
end 12'h41e:    begin Red = 8'hc2;    Green = 8'h9b;    Blue = 8'h6d;
end 12'h41f:    begin Red = 8'hb8;    Green = 8'h8a;    Blue = 8'h58;
end 12'h420:    begin Red = 8'hb4;    Green = 8'h87;    Blue = 8'h62;
end 12'h421:    begin Red = 8'h79;    Green = 8'h87;    Blue = 8'h10;
end 12'h422:    begin Red = 8'h80;    Green = 8'h88;    Blue = 8'h19;
end 12'h423:    begin Red = 8'h63;    Green = 8'h51;    Blue = 8'h23;
end 12'h424:    begin Red = 8'h4f;    Green = 8'h44;    Blue = 8'h2b;
end 12'h425:    begin Red = 8'h0a;    Green = 8'h0b;    Blue = 8'hbb;
end 12'h426:    begin Red = 8'h0a;    Green = 8'h4b;    Blue = 8'hae;
end 12'h427:    begin Red = 8'h09;    Green = 8'hdb;    Blue = 8'h9d;
end 12'h428:    begin Red = 8'h6f;    Green = 8'h7b;    Blue = 8'h21;
end 12'h429:    begin Red = 8'h08;    Green = 8'hba;    Blue = 8'h79;
end 12'h42a:    begin Red = 8'h48;    Green = 8'h37;    Blue = 8'h1d;
end 12'h42b:    begin Red = 8'h40;    Green = 8'h3e;    Blue = 8'h1f;
end 12'h42c:    begin Red = 8'h4d;    Green = 8'h42;    Blue = 8'h1e;
end 12'h42d:    begin Red = 8'hbd;    Green = 8'h9a;    Blue = 8'h79;
end 12'h42e:    begin Red = 8'h07;    Green = 8'hb7;    Blue = 8'hee;
end 12'h42f:    begin Red = 8'h66;    Green = 8'h63;    Blue = 8'h31;
end 12'h430:    begin Red = 8'h84;    Green = 8'h7f;    Blue = 8'h26;
end 12'h431:    begin Red = 8'hbc;    Green = 8'hae;    Blue = 8'h36;
end 12'h432:    begin Red = 8'h84;    Green = 8'h84;    Blue = 8'h26;
end 12'h433:    begin Red = 8'h92;    Green = 8'h87;    Blue = 8'h2d;
end 12'h434:    begin Red = 8'h86;    Green = 8'h6a;    Blue = 8'h55;
end 12'h435:    begin Red = 8'h7e;    Green = 8'h62;    Blue = 8'h4d;
end 12'h436:    begin Red = 8'h9d;    Green = 8'h8a;    Blue = 8'h5e;
end 12'h437:    begin Red = 8'haf;    Green = 8'hb0;    Blue = 8'hb5;
end 12'h438:    begin Red = 8'hc7;    Green = 8'hc6;    Blue = 8'hc5;
end 12'h439:    begin Red = 8'h6b;    Green = 8'h71;    Blue = 8'h24;
end 12'h43a:    begin Red = 8'h6f;    Green = 8'h70;    Blue = 8'h2d;
end 12'h43b:    begin Red = 8'h7e;    Green = 8'h9d;    Blue = 8'h29;
end 12'h43c:    begin Red = 8'hbb;    Green = 8'h8f;    Blue = 8'h5c;
end 12'h43d:    begin Red = 8'hbb;    Green = 8'h93;    Blue = 8'h61;
end 12'h43e:    begin Red = 8'h80;    Green = 8'h87;    Blue = 8'h13;
end 12'h43f:    begin Red = 8'h59;    Green = 8'h5f;    Blue = 8'h2b;
end 12'h440:    begin Red = 8'h40;    Green = 8'h3d;    Blue = 8'h2d;
end 12'h441:    begin Red = 8'h6b;    Green = 8'h63;    Blue = 8'h34;
end 12'h442:    begin Red = 8'h4c;    Green = 8'h45;    Blue = 8'h25;
end 12'h443:    begin Red = 8'h91;    Green = 8'hac;    Blue = 8'h15;
end 12'h444:    begin Red = 8'h3b;    Green = 8'h30;    Blue = 8'h24;
end 12'h445:    begin Red = 8'h3e;    Green = 8'h2e;    Blue = 8'h29;
end 12'h446:    begin Red = 8'h02;    Green = 8'h53;    Blue = 8'h5c;
end 12'h447:    begin Red = 8'h9f;    Green = 8'h87;    Blue = 8'h59;
end 12'h448:    begin Red = 8'h9f;    Green = 8'hc9;    Blue = 8'h1b;
end 12'h449:    begin Red = 8'h93;    Green = 8'hb4;    Blue = 8'h23;
end 12'h44a:    begin Red = 8'ha6;    Green = 8'hc4;    Blue = 8'h18;
end 12'h44b:    begin Red = 8'h95;    Green = 8'h78;    Blue = 8'h51;
end 12'h44c:    begin Red = 8'hb7;    Green = 8'hb2;    Blue = 8'h1a;
end 12'h44d:    begin Red = 8'h8a;    Green = 8'h8d;    Blue = 8'h9d;
end 12'h44e:    begin Red = 8'h91;    Green = 8'h90;    Blue = 8'h91;
end 12'h44f:    begin Red = 8'h69;    Green = 8'h81;    Blue = 8'h7b;
end 12'h450:    begin Red = 8'h49;    Green = 8'h5f;    Blue = 8'h11;
end 12'h451:    begin Red = 8'h5b;    Green = 8'h74;    Blue = 8'h66;
end 12'h452:    begin Red = 8'h57;    Green = 8'h79;    Blue = 8'h5f;
end 12'h453:    begin Red = 8'hd8;    Green = 8'ha9;    Blue = 8'h7d;
end 12'h454:    begin Red = 8'h8d;    Green = 8'h90;    Blue = 8'h19;
end 12'h455:    begin Red = 8'h09;    Green = 8'h2b;    Blue = 8'h6b;
end 12'h456:    begin Red = 8'h6a;    Green = 8'h81;    Blue = 8'h32;
end 12'h457:    begin Red = 8'h3f;    Green = 8'h3c;    Blue = 8'h27;
end 12'h458:    begin Red = 8'ha4;    Green = 8'hce;    Blue = 8'h22;
end 12'h459:    begin Red = 8'h41;    Green = 8'h38;    Blue = 8'h2c;
end 12'h45a:    begin Red = 8'h08;    Green = 8'hca;    Blue = 8'hfb;
end 12'h45b:    begin Red = 8'h09;    Green = 8'h1b;    Blue = 8'hcc;
end 12'h45c:    begin Red = 8'h37;    Green = 8'h2f;    Blue = 8'h1f;
end 12'h45d:    begin Red = 8'h08;    Green = 8'hcb;    Blue = 8'h26;
end 12'h45e:    begin Red = 8'h3a;    Green = 8'h29;    Blue = 8'h2d;
end 12'h45f:    begin Red = 8'hbf;    Green = 8'h9e;    Blue = 8'h86;
end 12'h460:    begin Red = 8'h07;    Green = 8'hc7;    Blue = 8'h58;
end 12'h461:    begin Red = 8'h85;    Green = 8'h81;    Blue = 8'h20;
end 12'h462:    begin Red = 8'h0a;    Green = 8'hdd;    Blue = 8'h6d;
end 12'h463:    begin Red = 8'h44;    Green = 8'h38;    Blue = 8'h3d;
end 12'h464:    begin Red = 8'h08;    Green = 8'hfa;    Blue = 8'hcb;
end 12'h465:    begin Red = 8'h5a;    Green = 8'h63;    Blue = 8'h3d;
end 12'h466:    begin Red = 8'h59;    Green = 8'h63;    Blue = 8'h38;
end 12'h467:    begin Red = 8'h97;    Green = 8'h7d;    Blue = 8'h44;
end 12'h468:    begin Red = 8'h08;    Green = 8'hf8;    Blue = 8'hef;
end 12'h469:    begin Red = 8'hbc;    Green = 8'hb3;    Blue = 8'h2e;
end 12'h46a:    begin Red = 8'hbf;    Green = 8'hbd;    Blue = 8'h20;
end 12'h46b:    begin Red = 8'h6b;    Green = 8'h51;    Blue = 8'h3c;
end 12'h46c:    begin Red = 8'h46;    Green = 8'h51;    Blue = 8'h23;
end 12'h46d:    begin Red = 8'h67;    Green = 8'h84;    Blue = 8'h65;
end 12'h46e:    begin Red = 8'h68;    Green = 8'h81;    Blue = 8'h73;
end 12'h46f:    begin Red = 8'h6c;    Green = 8'h84;    Blue = 8'h6e;
end 12'h470:    begin Red = 8'h5b;    Green = 8'h78;    Blue = 8'h18;
end 12'h471:    begin Red = 8'h83;    Green = 8'h95;    Blue = 8'h23;
end 12'h472:    begin Red = 8'h79;    Green = 8'h7f;    Blue = 8'h17;
end 12'h473:    begin Red = 8'h8d;    Green = 8'h89;    Blue = 8'h32;
end 12'h474:    begin Red = 8'h93;    Green = 8'h91;    Blue = 8'h22;
end 12'h475:    begin Red = 8'h58;    Green = 8'h56;    Blue = 8'h37;
end 12'h476:    begin Red = 8'h9a;    Green = 8'hc9;    Blue = 8'h19;
end 12'h477:    begin Red = 8'h09;    Green = 8'hdb;    Blue = 8'hcd;
end 12'h478:    begin Red = 8'h08;    Green = 8'h9a;    Blue = 8'h5b;
end 12'h479:    begin Red = 8'h08;    Green = 8'haa;    Blue = 8'h5e;
end 12'h47a:    begin Red = 8'he0;    Green = 8'ha5;    Blue = 8'h76;
end 12'h47b:    begin Red = 8'h4b;    Green = 8'h4f;    Blue = 8'h26;
end 12'h47c:    begin Red = 8'h87;    Green = 8'h87;    Blue = 8'h10;
end 12'h47d:    begin Red = 8'h44;    Green = 8'h38;    Blue = 8'h24;
end 12'h47e:    begin Red = 8'h6d;    Green = 8'h66;    Blue = 8'h2a;
end 12'h47f:    begin Red = 8'h69;    Green = 8'h5d;    Blue = 8'h25;
end 12'h480:    begin Red = 8'h02;    Green = 8'h43;    Blue = 8'h5e;
end 12'h481:    begin Red = 8'h84;    Green = 8'h65;    Blue = 8'h49;
end 12'h482:    begin Red = 8'ha0;    Green = 8'h85;    Blue = 8'h6b;
end 12'h483:    begin Red = 8'hb8;    Green = 8'h94;    Blue = 8'h76;
end 12'h484:    begin Red = 8'h0a;    Green = 8'h7a;    Blue = 8'h12;
end 12'h485:    begin Red = 8'h90;    Green = 8'h7f;    Blue = 8'h49;
end 12'h486:    begin Red = 8'hbb;    Green = 8'ha3;    Blue = 8'h70;
end 12'h487:    begin Red = 8'h08;    Green = 8'h68;    Blue = 8'hed;
end 12'h488:    begin Red = 8'h90;    Green = 8'h7d;    Blue = 8'h53;
end 12'h489:    begin Red = 8'hb8;    Green = 8'h9b;    Blue = 8'h6c;
end 12'h48a:    begin Red = 8'hd6;    Green = 8'h98;    Blue = 8'h64;
end 12'h48b:    begin Red = 8'ha5;    Green = 8'hb0;    Blue = 8'h19;
end 12'h48c:    begin Red = 8'h63;    Green = 8'h6f;    Blue = 8'h38;
end 12'h48d:    begin Red = 8'h08;    Green = 8'h29;    Blue = 8'hbf;
end 12'h48e:    begin Red = 8'h02;    Green = 8'h42;    Blue = 8'h6e;
end 12'h48f:    begin Red = 8'h9f;    Green = 8'h77;    Blue = 8'h4a;
end 12'h490:    begin Red = 8'h03;    Green = 8'hd2;    Blue = 8'hd9;
end 12'h491:    begin Red = 8'h47;    Green = 8'h33;    Blue = 8'h15;
end 12'h492:    begin Red = 8'h6a;    Green = 8'h5d;    Blue = 8'h2b;
end 12'h493:    begin Red = 8'h03;    Green = 8'hc3;    Blue = 8'h1e;
end 12'h494:    begin Red = 8'h36;    Green = 8'h30;    Blue = 8'h13;
end 12'h495:    begin Red = 8'h52;    Green = 8'h53;    Blue = 8'h22;
end 12'h496:    begin Red = 8'h08;    Green = 8'h7a;    Blue = 8'h2a;
end 12'h497:    begin Red = 8'h21;    Green = 8'h25;    Blue = 8'h15;
end 12'h498:    begin Red = 8'h9d;    Green = 8'h81;    Blue = 8'h52;
end 12'h499:    begin Red = 8'he2;    Green = 8'hc8;    Blue = 8'h95;
end 12'h49a:    begin Red = 8'he6;    Green = 8'hc5;    Blue = 8'ha5;
end 12'h49b:    begin Red = 8'h8e;    Green = 8'h7a;    Blue = 8'h3e;
end 12'h49c:    begin Red = 8'he0;    Green = 8'hc7;    Blue = 8'h81;
end 12'h49d:    begin Red = 8'h80;    Green = 8'h87;    Blue = 8'h90;
end 12'h49e:    begin Red = 8'h8a;    Green = 8'h8d;    Blue = 8'h8d;
end 12'h49f:    begin Red = 8'ha6;    Green = 8'ha9;    Blue = 8'ha8;
end 12'h4a0:    begin Red = 8'hab;    Green = 8'haa;    Blue = 8'hab;
end 12'h4a1:    begin Red = 8'h02;    Green = 8'h92;    Blue = 8'hfe;
end 12'h4a2:    begin Red = 8'h88;    Green = 8'h9a;    Blue = 8'h15;
end 12'h4a3:    begin Red = 8'h81;    Green = 8'h95;    Blue = 8'h18;
end 12'h4a4:    begin Red = 8'h9b;    Green = 8'hab;    Blue = 8'h22;
end 12'h4a5:    begin Red = 8'h02;    Green = 8'he3;    Blue = 8'h8e;
end 12'h4a6:    begin Red = 8'h01;    Green = 8'h02;    Blue = 8'h60;
end 12'h4a7:    begin Red = 8'h02;    Green = 8'h72;    Blue = 8'hae;
end 12'h4a8:    begin Red = 8'hba;    Green = 8'h84;    Blue = 8'h4c;
end 12'h4a9:    begin Red = 8'h02;    Green = 8'h22;    Blue = 8'h79;
end 12'h4aa:    begin Red = 8'h02;    Green = 8'h82;    Blue = 8'h3e;
end 12'h4ab:    begin Red = 8'h53;    Green = 8'h53;    Blue = 8'h27;
end 12'h4ac:    begin Red = 8'ha7;    Green = 8'h7f;    Blue = 8'h43;
end 12'h4ad:    begin Red = 8'h5f;    Green = 8'h58;    Blue = 8'h28;
end 12'h4ae:    begin Red = 8'h03;    Green = 8'hd3;    Blue = 8'h7e;
end 12'h4af:    begin Red = 8'h02;    Green = 8'he3;    Blue = 8'h9c;
end 12'h4b0:    begin Red = 8'h02;    Green = 8'h12;    Blue = 8'hd3;
end 12'h4b1:    begin Red = 8'h74;    Green = 8'h85;    Blue = 8'h2e;
end 12'h4b2:    begin Red = 8'h7a;    Green = 8'h5f;    Blue = 8'h3b;
end 12'h4b3:    begin Red = 8'hcc;    Green = 8'haf;    Blue = 8'h7e;
end 12'h4b4:    begin Red = 8'hc7;    Green = 8'hc3;    Blue = 8'h1a;
end 12'h4b5:    begin Red = 8'h82;    Green = 8'h7c;    Blue = 8'h37;
end 12'h4b6:    begin Red = 8'h02;    Green = 8'h32;    Blue = 8'hce;
end 12'h4b7:    begin Red = 8'hab;    Green = 8'h80;    Blue = 8'h65;
end 12'h4b8:    begin Red = 8'hff;    Green = 8'hd8;    Blue = 8'ha9;
end 12'h4b9:    begin Red = 8'hee;    Green = 8'hc5;    Blue = 8'h97;
end 12'h4ba:    begin Red = 8'he8;    Green = 8'hc4;    Blue = 8'h94;
end 12'h4bb:    begin Red = 8'he9;    Green = 8'hcc;    Blue = 8'h9e;
end 12'h4bc:    begin Red = 8'h7a;    Green = 8'h83;    Blue = 8'h89;
end 12'h4bd:    begin Red = 8'hdd;    Green = 8'hb2;    Blue = 8'h83;
end 12'h4be:    begin Red = 8'hd4;    Green = 8'ha2;    Blue = 8'h6f;
end 12'h4bf:    begin Red = 8'hbb;    Green = 8'hb5;    Blue = 8'h21;
end 12'h4c0:    begin Red = 8'h81;    Green = 8'h7d;    Blue = 8'h2d;
end 12'h4c1:    begin Red = 8'ha1;    Green = 8'hbc;    Blue = 8'h23;
end 12'h4c2:    begin Red = 8'h01;    Green = 8'h02;    Blue = 8'h50;
end 12'h4c3:    begin Red = 8'he7;    Green = 8'haa;    Blue = 8'h7c;
end 12'h4c4:    begin Red = 8'hee;    Green = 8'hac;    Blue = 8'h7c;
end 12'h4c5:    begin Red = 8'h3c;    Green = 8'h35;    Blue = 8'h11;
end 12'h4c6:    begin Red = 8'h45;    Green = 8'h2f;    Blue = 8'h10;
end 12'h4c7:    begin Red = 8'h9d;    Green = 8'h71;    Blue = 8'h3d;
end 12'h4c8:    begin Red = 8'hb1;    Green = 8'h7b;    Blue = 8'h4f;
end 12'h4c9:    begin Red = 8'ha7;    Green = 8'h77;    Blue = 8'h40;
end 12'h4ca:    begin Red = 8'ha7;    Green = 8'h7a;    Blue = 8'h48;
end 12'h4cb:    begin Red = 8'hb5;    Green = 8'h74;    Blue = 8'h56;
end 12'h4cc:    begin Red = 8'ha5;    Green = 8'h70;    Blue = 8'h48;
end 12'h4cd:    begin Red = 8'h04;    Green = 8'h13;    Blue = 8'hab;
end 12'h4ce:    begin Red = 8'h3d;    Green = 8'h30;    Blue = 8'h16;
end 12'h4cf:    begin Red = 8'h02;    Green = 8'hc2;    Blue = 8'h8b;
end 12'h4d0:    begin Red = 8'h8c;    Green = 8'h70;    Blue = 8'h44;
end 12'h4d1:    begin Red = 8'h08;    Green = 8'h09;    Blue = 8'h9f;
end 12'h4d2:    begin Red = 8'hb0;    Green = 8'hcf;    Blue = 8'h1f;
end 12'h4d3:    begin Red = 8'ha2;    Green = 8'ha8;    Blue = 8'haf;
end 12'h4d4:    begin Red = 8'hc2;    Green = 8'h77;    Blue = 8'haf;
end 12'h4d5:    begin Red = 8'hc5;    Green = 8'h7a;    Blue = 8'h9b;
end 12'h4d6:    begin Red = 8'hbc;    Green = 8'h7f;    Blue = 8'had;
end 12'h4d7:    begin Red = 8'hca;    Green = 8'hd7;    Blue = 8'hcb;
end 12'h4d8:    begin Red = 8'hd0;    Green = 8'hbe;    Blue = 8'h99;
end 12'h4d9:    begin Red = 8'h02;    Green = 8'hd3;    Blue = 8'h4e;
end 12'h4da:    begin Red = 8'h08;    Green = 8'h1a;    Blue = 8'h1e;
end 12'h4db:    begin Red = 8'hb6;    Green = 8'h94;    Blue = 8'h5a;
end 12'h4dc:    begin Red = 8'h95;    Green = 8'h80;    Blue = 8'h29;
end 12'h4dd:    begin Red = 8'hbd;    Green = 8'hb2;    Blue = 8'h26;
end 12'h4de:    begin Red = 8'h5f;    Green = 8'h63;    Blue = 8'h2b;
end 12'h4df:    begin Red = 8'h08;    Green = 8'h8a;    Blue = 8'h3d;
end 12'h4e0:    begin Red = 8'h09;    Green = 8'h0a;    Blue = 8'hce;
end 12'h4e1:    begin Red = 8'h66;    Green = 8'h56;    Blue = 8'h1f;
end 12'h4e2:    begin Red = 8'h2c;    Green = 8'h2a;    Blue = 8'h10;
end 12'h4e3:    begin Red = 8'hab;    Green = 8'h83;    Blue = 8'h48;
end 12'h4e4:    begin Red = 8'hc6;    Green = 8'h7e;    Blue = 8'h52;
end 12'h4e5:    begin Red = 8'h35;    Green = 8'h29;    Blue = 8'h10;
end 12'h4e6:    begin Red = 8'h3a;    Green = 8'h25;    Blue = 8'h11;
end 12'h4e7:    begin Red = 8'h02;    Green = 8'h82;    Blue = 8'hcb;
end 12'h4e8:    begin Red = 8'h6d;    Green = 8'h5c;    Blue = 8'h1e;
end 12'h4e9:    begin Red = 8'h6d;    Green = 8'h5d;    Blue = 8'h18;
end 12'h4ea:    begin Red = 8'h6c;    Green = 8'h56;    Blue = 8'h17;
end 12'h4eb:    begin Red = 8'h04;    Green = 8'hf4;    Blue = 8'hdd;
end 12'h4ec:    begin Red = 8'hff;    Green = 8'hd9;    Blue = 8'hb0;
end 12'h4ed:    begin Red = 8'h5c;    Green = 8'h40;    Blue = 8'h38;
end 12'h4ee:    begin Red = 8'hd0;    Green = 8'haf;    Blue = 8'h90;
end 12'h4ef:    begin Red = 8'hd7;    Green = 8'hb4;    Blue = 8'ha9;
end 12'h4f0:    begin Red = 8'hce;    Green = 8'ha4;    Blue = 8'hab;
end 12'h4f1:    begin Red = 8'hc1;    Green = 8'hb1;    Blue = 8'h36;
end 12'h4f2:    begin Red = 8'h81;    Green = 8'h77;    Blue = 8'h1c;
end 12'h4f3:    begin Red = 8'hcc;    Green = 8'hba;    Blue = 8'h33;
end 12'h4f4:    begin Red = 8'ha4;    Green = 8'h96;    Blue = 8'h27;
end 12'h4f5:    begin Red = 8'h52;    Green = 8'h4c;    Blue = 8'h37;
end 12'h4f6:    begin Red = 8'h96;    Green = 8'hb9;    Blue = 8'h12;
end 12'h4f7:    begin Red = 8'h2c;    Green = 8'h1a;    Blue = 8'h32;
end 12'h4f8:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'hfa;
end 12'h4f9:    begin Red = 8'hf7;    Green = 8'hc8;    Blue = 8'h9e;
end 12'h4fa:    begin Red = 8'had;    Green = 8'h55;    Blue = 8'h95;
end 12'h4fb:    begin Red = 8'ha3;    Green = 8'h52;    Blue = 8'h95;
end 12'h4fc:    begin Red = 8'hc6;    Green = 8'hd8;    Blue = 8'hd9;
end 12'h4fd:    begin Red = 8'hc5;    Green = 8'hda;    Blue = 8'hcb;
end 12'h4fe:    begin Red = 8'hc6;    Green = 8'hcd;    Blue = 8'hc3;
end 12'h4ff:    begin Red = 8'hf1;    Green = 8'he5;    Blue = 8'hc0;
end 12'h500:    begin Red = 8'hf0;    Green = 8'he6;    Blue = 8'hb7;
end 12'h501:    begin Red = 8'hcc;    Green = 8'hc1;    Blue = 8'h93;
end 12'h502:    begin Red = 8'hcf;    Green = 8'hcc;    Blue = 8'h93;
end 12'h503:    begin Red = 8'h95;    Green = 8'hae;    Blue = 8'h88;
end 12'h504:    begin Red = 8'h5c;    Green = 8'h7f;    Blue = 8'h61;
end 12'h505:    begin Red = 8'h48;    Green = 8'h48;    Blue = 8'h42;
end 12'h506:    begin Red = 8'h66;    Green = 8'h75;    Blue = 8'h72;
end 12'h507:    begin Red = 8'h5c;    Green = 8'h71;    Blue = 8'h6c;
end 12'h508:    begin Red = 8'h4d;    Green = 8'h6f;    Blue = 8'h66;
end 12'h509:    begin Red = 8'hdd;    Green = 8'h9f;    Blue = 8'h78;
end 12'h50a:    begin Red = 8'hc8;    Green = 8'haf;    Blue = 8'h2f;
end 12'h50b:    begin Red = 8'h85;    Green = 8'h7a;    Blue = 8'h21;
end 12'h50c:    begin Red = 8'h8f;    Green = 8'h83;    Blue = 8'h32;
end 12'h50d:    begin Red = 8'h61;    Green = 8'h6c;    Blue = 8'h3d;
end 12'h50e:    begin Red = 8'h00;    Green = 8'hcf;    Blue = 8'h13;
end 12'h50f:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'hee;
end 12'h510:    begin Red = 8'h03;    Green = 8'h53;    Blue = 8'hd9;
end 12'h511:    begin Red = 8'h02;    Green = 8'ha3;    Blue = 8'h4d;
end 12'h512:    begin Red = 8'h5f;    Green = 8'h55;    Blue = 8'h1e;
end 12'h513:    begin Red = 8'h03;    Green = 8'hf3;    Blue = 8'h6f;
end 12'h514:    begin Red = 8'hb7;    Green = 8'h81;    Blue = 8'h55;
end 12'h515:    begin Red = 8'h72;    Green = 8'h68;    Blue = 8'h30;
end 12'h516:    begin Red = 8'h03;    Green = 8'he3;    Blue = 8'h5e;
end 12'h517:    begin Red = 8'h42;    Green = 8'h34;    Blue = 8'h12;
end 12'h518:    begin Red = 8'h6c;    Green = 8'h4f;    Blue = 8'h1d;
end 12'h519:    begin Red = 8'h61;    Green = 8'h50;    Blue = 8'h1c;
end 12'h51a:    begin Red = 8'hee;    Green = 8'hc8;    Blue = 8'ha4;
end 12'h51b:    begin Red = 8'h6c;    Green = 8'h77;    Blue = 8'h38;
end 12'h51c:    begin Red = 8'hb1;    Green = 8'h87;    Blue = 8'h7b;
end 12'h51d:    begin Red = 8'hac;    Green = 8'h86;    Blue = 8'h68;
end 12'h51e:    begin Red = 8'h7d;    Green = 8'h6c;    Blue = 8'h53;
end 12'h51f:    begin Red = 8'hc1;    Green = 8'h9f;    Blue = 8'h8d;
end 12'h520:    begin Red = 8'hb3;    Green = 8'hae;    Blue = 8'h2b;
end 12'h521:    begin Red = 8'h9f;    Green = 8'haf;    Blue = 8'h28;
end 12'h522:    begin Red = 8'h73;    Green = 8'h77;    Blue = 8'h36;
end 12'h523:    begin Red = 8'hff;    Green = 8'hc7;    Blue = 8'hab;
end 12'h524:    begin Red = 8'hc5;    Green = 8'hac;    Blue = 8'h81;
end 12'h525:    begin Red = 8'haf;    Green = 8'h6a;    Blue = 8'h99;
end 12'h526:    begin Red = 8'hbf;    Green = 8'hc5;    Blue = 8'hc3;
end 12'h527:    begin Red = 8'h82;    Green = 8'h9d;    Blue = 8'h6d;
end 12'h528:    begin Red = 8'he9;    Green = 8'he1;    Blue = 8'hb6;
end 12'h529:    begin Red = 8'h84;    Green = 8'h99;    Blue = 8'h7a;
end 12'h52a:    begin Red = 8'h02;    Green = 8'h52;    Blue = 8'hec;
end 12'h52b:    begin Red = 8'h63;    Green = 8'h7e;    Blue = 8'h6d;
end 12'h52c:    begin Red = 8'h80;    Green = 8'h7e;    Blue = 8'h21;
end 12'h52d:    begin Red = 8'hbc;    Green = 8'hac;    Blue = 8'h3f;
end 12'h52e:    begin Red = 8'h68;    Green = 8'h5d;    Blue = 8'h38;
end 12'h52f:    begin Red = 8'had;    Green = 8'hca;    Blue = 8'h18;
end 12'h530:    begin Red = 8'h94;    Green = 8'ha9;    Blue = 8'h1b;
end 12'h531:    begin Red = 8'h09;    Green = 8'h8c;    Blue = 8'h06;
end 12'h532:    begin Red = 8'h99;    Green = 8'hb3;    Blue = 8'h12;
end 12'h533:    begin Red = 8'h01;    Green = 8'hc1;    Blue = 8'hfc;
end 12'h534:    begin Red = 8'h03;    Green = 8'h03;    Blue = 8'h8e;
end 12'h535:    begin Red = 8'h9c;    Green = 8'h76;    Blue = 8'h41;
end 12'h536:    begin Red = 8'h03;    Green = 8'hb3;    Blue = 8'h2e;
end 12'h537:    begin Red = 8'h67;    Green = 8'h50;    Blue = 8'h16;
end 12'h538:    begin Red = 8'h03;    Green = 8'hd3;    Blue = 8'h0b;
end 12'h539:    begin Red = 8'h5d;    Green = 8'h4b;    Blue = 8'h17;
end 12'h53a:    begin Red = 8'h07;    Green = 8'h67;    Blue = 8'h88;
end 12'h53b:    begin Red = 8'hb7;    Green = 8'hab;    Blue = 8'h30;
end 12'h53c:    begin Red = 8'h87;    Green = 8'hac;    Blue = 8'h16;
end 12'h53d:    begin Red = 8'h72;    Green = 8'h61;    Blue = 8'h3f;
end 12'h53e:    begin Red = 8'ha4;    Green = 8'h58;    Blue = 8'h8d;
end 12'h53f:    begin Red = 8'hbf;    Green = 8'h75;    Blue = 8'ha5;
end 12'h540:    begin Red = 8'hc5;    Green = 8'h80;    Blue = 8'hac;
end 12'h541:    begin Red = 8'he1;    Green = 8'hd7;    Blue = 8'hac;
end 12'h542:    begin Red = 8'h02;    Green = 8'h83;    Blue = 8'h10;
end 12'h543:    begin Red = 8'h65;    Green = 8'h63;    Blue = 8'h2a;
end 12'h544:    begin Red = 8'h47;    Green = 8'h44;    Blue = 8'h1d;
end 12'h545:    begin Red = 8'h4c;    Green = 8'h3f;    Blue = 8'h29;
end 12'h546:    begin Red = 8'haa;    Green = 8'hcc;    Blue = 8'h21;
end 12'h547:    begin Red = 8'h49;    Green = 8'h3d;    Blue = 8'h21;
end 12'h548:    begin Red = 8'h68;    Green = 8'h57;    Blue = 8'h24;
end 12'h549:    begin Red = 8'h96;    Green = 8'h67;    Blue = 8'h2b;
end 12'h54a:    begin Red = 8'h8a;    Green = 8'h62;    Blue = 8'h27;
end 12'h54b:    begin Red = 8'h03;    Green = 8'h62;    Blue = 8'hbd;
end 12'h54c:    begin Red = 8'h03;    Green = 8'h03;    Blue = 8'h0e;
end 12'h54d:    begin Red = 8'h89;    Green = 8'h56;    Blue = 8'h23;
end 12'h54e:    begin Red = 8'h82;    Green = 8'h54;    Blue = 8'h1d;
end 12'h54f:    begin Red = 8'h52;    Green = 8'h41;    Blue = 8'h30;
end 12'h550:    begin Red = 8'hcb;    Green = 8'hc2;    Blue = 8'h2c;
end 12'h551:    begin Red = 8'h86;    Green = 8'h89;    Blue = 8'h26;
end 12'h552:    begin Red = 8'he1;    Green = 8'hd0;    Blue = 8'h2d;
end 12'h553:    begin Red = 8'h03;    Green = 8'h62;    Blue = 8'hdf;
end 12'h554:    begin Red = 8'h33;    Green = 8'h19;    Blue = 8'h34;
end 12'h555:    begin Red = 8'h8a;    Green = 8'ha9;    Blue = 8'h1b;
end 12'h556:    begin Red = 8'h97;    Green = 8'hbb;    Blue = 8'h1b;
end 12'h557:    begin Red = 8'h72;    Green = 8'h64;    Blue = 8'h37;
end 12'h558:    begin Red = 8'h48;    Green = 8'h64;    Blue = 8'h10;
end 12'h559:    begin Red = 8'hb3;    Green = 8'h6d;    Blue = 8'ha1;
end 12'h55a:    begin Red = 8'hac;    Green = 8'h5b;    Blue = 8'h8c;
end 12'h55b:    begin Red = 8'hc7;    Green = 8'hd6;    Blue = 8'hbe;
end 12'h55c:    begin Red = 8'hc6;    Green = 8'he3;    Blue = 8'hca;
end 12'h55d:    begin Red = 8'hc1;    Green = 8'h86;    Blue = 8'hbd;
end 12'h55e:    begin Red = 8'hf5;    Green = 8'hed;    Blue = 8'hbf;
end 12'h55f:    begin Red = 8'h09;    Green = 8'hc8;    Blue = 8'hdc;
end 12'h560:    begin Red = 8'h8f;    Green = 8'h90;    Blue = 8'h10;
end 12'h561:    begin Red = 8'h74;    Green = 8'h87;    Blue = 8'h64;
end 12'h562:    begin Red = 8'h9c;    Green = 8'h7a;    Blue = 8'h57;
end 12'h563:    begin Red = 8'hb6;    Green = 8'hb4;    Blue = 8'h21;
end 12'h564:    begin Red = 8'h9e;    Green = 8'h87;    Blue = 8'h2b;
end 12'h565:    begin Red = 8'h89;    Green = 8'h8e;    Blue = 8'h25;
end 12'h566:    begin Red = 8'hc8;    Green = 8'hc0;    Blue = 8'h34;
end 12'h567:    begin Red = 8'h03;    Green = 8'h42;    Blue = 8'hbc;
end 12'h568:    begin Red = 8'hae;    Green = 8'hcd;    Blue = 8'h27;
end 12'h569:    begin Red = 8'h97;    Green = 8'h67;    Blue = 8'h30;
end 12'h56a:    begin Red = 8'h8a;    Green = 8'h66;    Blue = 8'h2d;
end 12'h56b:    begin Red = 8'h5e;    Green = 8'h51;    Blue = 8'h17;
end 12'h56c:    begin Red = 8'h85;    Green = 8'h4e;    Blue = 8'h20;
end 12'h56d:    begin Red = 8'h7f;    Green = 8'h52;    Blue = 8'h23;
end 12'h56e:    begin Red = 8'h8a;    Green = 8'h72;    Blue = 8'h3d;
end 12'h56f:    begin Red = 8'hcd;    Green = 8'hbc;    Blue = 8'h2d;
end 12'h570:    begin Red = 8'h49;    Green = 8'h59;    Blue = 8'h25;
end 12'h571:    begin Red = 8'hc0;    Green = 8'haa;    Blue = 8'h2d;
end 12'h572:    begin Red = 8'hd8;    Green = 8'hca;    Blue = 8'h36;
end 12'h573:    begin Red = 8'h08;    Green = 8'hba;    Blue = 8'hbf;
end 12'h574:    begin Red = 8'h5c;    Green = 8'h77;    Blue = 8'h23;
end 12'h575:    begin Red = 8'had;    Green = 8'h56;    Blue = 8'h9d;
end 12'h576:    begin Red = 8'hce;    Green = 8'hc4;    Blue = 8'hcc;
end 12'h577:    begin Red = 8'hc4;    Green = 8'hdd;    Blue = 8'hd3;
end 12'h578:    begin Red = 8'hd2;    Green = 8'hca;    Blue = 8'ha4;
end 12'h579:    begin Red = 8'hcc;    Green = 8'hc5;    Blue = 8'h98;
end 12'h57a:    begin Red = 8'hc1;    Green = 8'hc1;    Blue = 8'h8c;
end 12'h57b:    begin Red = 8'h9a;    Green = 8'h81;    Blue = 8'h2b;
end 12'h57c:    begin Red = 8'h53;    Green = 8'h53;    Blue = 8'h33;
end 12'h57d:    begin Red = 8'hb2;    Green = 8'haf;    Blue = 8'h20;
end 12'h57e:    begin Red = 8'ha7;    Green = 8'hc7;    Blue = 8'h11;
end 12'h57f:    begin Red = 8'ha5;    Green = 8'hcc;    Blue = 8'h11;
end 12'h580:    begin Red = 8'h08;    Green = 8'h8a;    Blue = 8'hbf;
end 12'h581:    begin Red = 8'h3c;    Green = 8'h4b;    Blue = 8'h27;
end 12'h582:    begin Red = 8'hba;    Green = 8'hb0;    Blue = 8'h89;
end 12'h583:    begin Red = 8'heb;    Green = 8'hd2;    Blue = 8'ha4;
end 12'h584:    begin Red = 8'h87;    Green = 8'h6f;    Blue = 8'h44;
end 12'h585:    begin Red = 8'hfc;    Green = 8'hdb;    Blue = 8'hc1;
end 12'h586:    begin Red = 8'hff;    Green = 8'hea;    Blue = 8'hd8;
end 12'h587:    begin Red = 8'h31;    Green = 8'h41;    Blue = 8'h1d;
end 12'h588:    begin Red = 8'h24;    Green = 8'h1a;    Blue = 8'h10;
end 12'h589:    begin Red = 8'h2e;    Green = 8'h20;    Blue = 8'h14;
end 12'h58a:    begin Red = 8'h71;    Green = 8'h62;    Blue = 8'h30;
end 12'h58b:    begin Red = 8'h36;    Green = 8'h2d;    Blue = 8'h25;
end 12'h58c:    begin Red = 8'h76;    Green = 8'h5e;    Blue = 8'h33;
end 12'h58d:    begin Red = 8'h71;    Green = 8'h61;    Blue = 8'h26;
end 12'h58e:    begin Red = 8'h3b;    Green = 8'h33;    Blue = 8'h29;
end 12'h58f:    begin Red = 8'h35;    Green = 8'h2f;    Blue = 8'h2b;
end 12'h590:    begin Red = 8'hb4;    Green = 8'hbd;    Blue = 8'hb3;
end 12'h591:    begin Red = 8'h9e;    Green = 8'hbd;    Blue = 8'h9d;
end 12'h592:    begin Red = 8'hcc;    Green = 8'h74;    Blue = 8'hb4;
end 12'h593:    begin Red = 8'hc2;    Green = 8'h70;    Blue = 8'ha6;
end 12'h594:    begin Red = 8'hef;    Green = 8'he0;    Blue = 8'ha8;
end 12'h595:    begin Red = 8'ha2;    Green = 8'hbc;    Blue = 8'h10;
end 12'h596:    begin Red = 8'h39;    Green = 8'h38;    Blue = 8'h2b;
end 12'h597:    begin Red = 8'h71;    Green = 8'h45;    Blue = 8'h3b;
end 12'h598:    begin Red = 8'h87;    Green = 8'h58;    Blue = 8'h49;
end 12'h599:    begin Red = 8'hc8;    Green = 8'hbb;    Blue = 8'h26;
end 12'h59a:    begin Red = 8'h25;    Green = 8'h3e;    Blue = 8'h11;
end 12'h59b:    begin Red = 8'h01;    Green = 8'hc1;    Blue = 8'hdd;
end 12'h59c:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h9e;
end 12'h59d:    begin Red = 8'h04;    Green = 8'h53;    Blue = 8'h7e;
end 12'h59e:    begin Red = 8'h40;    Green = 8'h2f;    Blue = 8'h22;
end 12'h59f:    begin Red = 8'h91;    Green = 8'h69;    Blue = 8'h31;
end 12'h5a0:    begin Red = 8'h85;    Green = 8'h61;    Blue = 8'h21;
end 12'h5a1:    begin Red = 8'h3a;    Green = 8'h3e;    Blue = 8'h20;
end 12'h5a2:    begin Red = 8'h9b;    Green = 8'h99;    Blue = 8'h73;
end 12'h5a3:    begin Red = 8'h62;    Green = 8'h4f;    Blue = 8'h2b;
end 12'h5a4:    begin Red = 8'h9c;    Green = 8'h82;    Blue = 8'h58;
end 12'h5a5:    begin Red = 8'hf0;    Green = 8'hd9;    Blue = 8'h9e;
end 12'h5a6:    begin Red = 8'h90;    Green = 8'h82;    Blue = 8'h22;
end 12'h5a7:    begin Red = 8'hac;    Green = 8'ha7;    Blue = 8'h25;
end 12'h5a8:    begin Red = 8'ha3;    Green = 8'h92;    Blue = 8'h2d;
end 12'h5a9:    begin Red = 8'h03;    Green = 8'he3;    Blue = 8'hae;
end 12'h5aa:    begin Red = 8'ha6;    Green = 8'hb0;    Blue = 8'h99;
end 12'h5ab:    begin Red = 8'hd0;    Green = 8'h84;    Blue = 8'hb7;
end 12'h5ac:    begin Red = 8'hcb;    Green = 8'h82;    Blue = 8'had;
end 12'h5ad:    begin Red = 8'hce;    Green = 8'h7c;    Blue = 8'hb2;
end 12'h5ae:    begin Red = 8'h5d;    Green = 8'h7d;    Blue = 8'h2d;
end 12'h5af:    begin Red = 8'h6c;    Green = 8'h66;    Blue = 8'h3f;
end 12'h5b0:    begin Red = 8'h78;    Green = 8'h57;    Blue = 8'h2d;
end 12'h5b1:    begin Red = 8'h89;    Green = 8'h5e;    Blue = 8'h33;
end 12'h5b2:    begin Red = 8'h03;    Green = 8'hc5;    Blue = 8'h0e;
end 12'h5b3:    begin Red = 8'h6a;    Green = 8'h52;    Blue = 8'h28;
end 12'h5b4:    begin Red = 8'h9d;    Green = 8'h69;    Blue = 8'h2a;
end 12'h5b5:    begin Red = 8'h8a;    Green = 8'h85;    Blue = 8'h5d;
end 12'h5b6:    begin Red = 8'h84;    Green = 8'h53;    Blue = 8'h22;
end 12'h5b7:    begin Red = 8'h58;    Green = 8'h45;    Blue = 8'h36;
end 12'h5b8:    begin Red = 8'hb7;    Green = 8'hb0;    Blue = 8'h32;
end 12'h5b9:    begin Red = 8'h4d;    Green = 8'h53;    Blue = 8'h1d;
end 12'h5ba:    begin Red = 8'h5e;    Green = 8'h52;    Blue = 8'h25;
end 12'h5bb:    begin Red = 8'h02;    Green = 8'hf2;    Blue = 8'heb;
end 12'h5bc:    begin Red = 8'h02;    Green = 8'h62;    Blue = 8'ha9;
end 12'h5bd:    begin Red = 8'h03;    Green = 8'h13;    Blue = 8'hcd;
end 12'h5be:    begin Red = 8'hd0;    Green = 8'hcb;    Blue = 8'hd1;
end 12'h5bf:    begin Red = 8'hc7;    Green = 8'hc1;    Blue = 8'h91;
end 12'h5c0:    begin Red = 8'h8a;    Green = 8'h89;    Blue = 8'h2b;
end 12'h5c1:    begin Red = 8'h8c;    Green = 8'ha7;    Blue = 8'h10;
end 12'h5c2:    begin Red = 8'h6a;    Green = 8'h7c;    Blue = 8'h75;
end 12'h5c3:    begin Red = 8'h4a;    Green = 8'h6f;    Blue = 8'h1a;
end 12'h5c4:    begin Red = 8'h40;    Green = 8'h30;    Blue = 8'h1b;
end 12'h5c5:    begin Red = 8'h46;    Green = 8'h39;    Blue = 8'h13;
end 12'h5c6:    begin Red = 8'hba;    Green = 8'h87;    Blue = 8'h52;
end 12'h5c7:    begin Red = 8'hee;    Green = 8'hea;    Blue = 8'hb1;
end 12'h5c8:    begin Red = 8'hc3;    Green = 8'hba;    Blue = 8'h9b;
end 12'h5c9:    begin Red = 8'h41;    Green = 8'h4c;    Blue = 8'h33;
end 12'h5ca:    begin Red = 8'h3f;    Green = 8'h48;    Blue = 8'h2e;
end 12'h5cb:    begin Red = 8'ha2;    Green = 8'h98;    Blue = 8'h71;
end 12'h5cc:    begin Red = 8'h8c;    Green = 8'h85;    Blue = 8'h63;
end 12'h5cd:    begin Red = 8'h8e;    Green = 8'h8b;    Blue = 8'h6a;
end 12'h5ce:    begin Red = 8'h87;    Green = 8'h72;    Blue = 8'h4f;
end 12'h5cf:    begin Red = 8'h5e;    Green = 8'h4f;    Blue = 8'h33;
end 12'h5d0:    begin Red = 8'h03;    Green = 8'ha5;    Blue = 8'hcb;
end 12'h5d1:    begin Red = 8'h53;    Green = 8'h76;    Blue = 8'h1c;
end 12'h5d2:    begin Red = 8'h03;    Green = 8'he3;    Blue = 8'h78;
end 12'h5d3:    begin Red = 8'hc3;    Green = 8'h86;    Blue = 8'h50;
end 12'h5d4:    begin Red = 8'hb3;    Green = 8'h84;    Blue = 8'h4e;
end 12'h5d5:    begin Red = 8'hbb;    Green = 8'h77;    Blue = 8'h48;
end 12'h5d6:    begin Red = 8'h03;    Green = 8'hc3;    Blue = 8'h7b;
end 12'h5d7:    begin Red = 8'hc8;    Green = 8'haa;    Blue = 8'h78;
end 12'h5d8:    begin Red = 8'h03;    Green = 8'hc4;    Blue = 8'h6e;
end 12'h5d9:    begin Red = 8'h66;    Green = 8'h7c;    Blue = 8'h2d;
end 12'h5da:    begin Red = 8'ha8;    Green = 8'hb1;    Blue = 8'hb1;
end 12'h5db:    begin Red = 8'hcd;    Green = 8'h79;    Blue = 8'hbb;
end 12'h5dc:    begin Red = 8'hc8;    Green = 8'h6e;    Blue = 8'hba;
end 12'h5dd:    begin Red = 8'hff;    Green = 8'hf6;    Blue = 8'hc6;
end 12'h5de:    begin Red = 8'hdd;    Green = 8'hcf;    Blue = 8'ha1;
end 12'h5df:    begin Red = 8'h57;    Green = 8'h6a;    Blue = 8'h4f;
end 12'h5e0:    begin Red = 8'h5b;    Green = 8'h6d;    Blue = 8'h58;
end 12'h5e1:    begin Red = 8'h83;    Green = 8'ha8;    Blue = 8'h8a;
end 12'h5e2:    begin Red = 8'h78;    Green = 8'ha5;    Blue = 8'h8e;
end 12'h5e3:    begin Red = 8'ha4;    Green = 8'hcb;    Blue = 8'h16;
end 12'h5e4:    begin Red = 8'h9c;    Green = 8'hc0;    Blue = 8'h14;
end 12'h5e5:    begin Red = 8'h3d;    Green = 8'h61;    Blue = 8'h11;
end 12'h5e6:    begin Red = 8'h3c;    Green = 8'h30;    Blue = 8'h10;
end 12'h5e7:    begin Red = 8'h02;    Green = 8'h72;    Blue = 8'h7b;
end 12'h5e8:    begin Red = 8'h01;    Green = 8'he2;    Blue = 8'h0b;
end 12'h5e9:    begin Red = 8'haf;    Green = 8'h76;    Blue = 8'h44;
end 12'h5ea:    begin Red = 8'h64;    Green = 8'h56;    Blue = 8'h32;
end 12'h5eb:    begin Red = 8'hf5;    Green = 8'hb2;    Blue = 8'h76;
end 12'h5ec:    begin Red = 8'hfa;    Green = 8'hbd;    Blue = 8'h82;
end 12'h5ed:    begin Red = 8'h4f;    Green = 8'h4c;    Blue = 8'h11;
end 12'h5ee:    begin Red = 8'hdd;    Green = 8'hd1;    Blue = 8'h99;
end 12'h5ef:    begin Red = 8'hb4;    Green = 8'ha9;    Blue = 8'h7e;
end 12'h5f0:    begin Red = 8'h84;    Green = 8'h62;    Blue = 8'h2c;
end 12'h5f1:    begin Red = 8'h62;    Green = 8'h56;    Blue = 8'h16;
end 12'h5f2:    begin Red = 8'h80;    Green = 8'h6a;    Blue = 8'h4b;
end 12'h5f3:    begin Red = 8'h4e;    Green = 8'h65;    Blue = 8'h11;
end 12'h5f4:    begin Red = 8'h03;    Green = 8'hf3;    Blue = 8'h2b;
end 12'h5f5:    begin Red = 8'h98;    Green = 8'h75;    Blue = 8'h46;
end 12'h5f6:    begin Red = 8'h5b;    Green = 8'h59;    Blue = 8'h23;
end 12'h5f7:    begin Red = 8'h03;    Green = 8'h44;    Blue = 8'h8f;
end 12'h5f8:    begin Red = 8'h71;    Green = 8'h7a;    Blue = 8'h30;
end 12'h5f9:    begin Red = 8'hc6;    Green = 8'h86;    Blue = 8'hc7;
end 12'h5fa:    begin Red = 8'hd1;    Green = 8'h71;    Blue = 8'ha6;
end 12'h5fb:    begin Red = 8'ha1;    Green = 8'hc3;    Blue = 8'h1a;
end 12'h5fc:    begin Red = 8'h5f;    Green = 8'h71;    Blue = 8'h7c;
end 12'h5fd:    begin Red = 8'h03;    Green = 8'h22;    Blue = 8'hfa;
end 12'h5fe:    begin Red = 8'h02;    Green = 8'h82;    Blue = 8'h36;
end 12'h5ff:    begin Red = 8'ha2;    Green = 8'h76;    Blue = 8'h3e;
end 12'h600:    begin Red = 8'h02;    Green = 8'h62;    Blue = 8'hcf;
end 12'h601:    begin Red = 8'he2;    Green = 8'hda;    Blue = 8'h9d;
end 12'h602:    begin Red = 8'hb7;    Green = 8'ha8;    Blue = 8'h83;
end 12'h603:    begin Red = 8'h83;    Green = 8'h8c;    Blue = 8'h4f;
end 12'h604:    begin Red = 8'h76;    Green = 8'h80;    Blue = 8'h53;
end 12'h605:    begin Red = 8'h71;    Green = 8'h78;    Blue = 8'h46;
end 12'h606:    begin Red = 8'h7c;    Green = 8'h4a;    Blue = 8'h10;
end 12'h607:    begin Red = 8'h7f;    Green = 8'h4b;    Blue = 8'h1c;
end 12'h608:    begin Red = 8'hee;    Green = 8'hc9;    Blue = 8'h9e;
end 12'h609:    begin Red = 8'h03;    Green = 8'ha3;    Blue = 8'h6e;
end 12'h60a:    begin Red = 8'h3b;    Green = 8'h35;    Blue = 8'h1f;
end 12'h60b:    begin Red = 8'h5e;    Green = 8'h52;    Blue = 8'h10;
end 12'h60c:    begin Red = 8'hb6;    Green = 8'ha7;    Blue = 8'hb7;
end 12'h60d:    begin Red = 8'hb5;    Green = 8'h62;    Blue = 8'h9c;
end 12'h60e:    begin Red = 8'hcd;    Green = 8'hd6;    Blue = 8'hc3;
end 12'h60f:    begin Red = 8'h87;    Green = 8'ha0;    Blue = 8'h6b;
end 12'h610:    begin Red = 8'h6d;    Green = 8'ha0;    Blue = 8'h8d;
end 12'h611:    begin Red = 8'h0a;    Green = 8'h0b;    Blue = 8'hff;
end 12'h612:    begin Red = 8'h03;    Green = 8'h12;    Blue = 8'hdf;
end 12'h613:    begin Red = 8'h03;    Green = 8'hf3;    Blue = 8'h85;
end 12'h614:    begin Red = 8'h04;    Green = 8'hd3;    Blue = 8'had;
end 12'h615:    begin Red = 8'hcb;    Green = 8'h9d;    Blue = 8'h5f;
end 12'h616:    begin Red = 8'h84;    Green = 8'h87;    Blue = 8'h53;
end 12'h617:    begin Red = 8'h3c;    Green = 8'h41;    Blue = 8'h25;
end 12'h618:    begin Red = 8'h06;    Green = 8'hd3;    Blue = 8'h40;
end 12'h619:    begin Red = 8'h06;    Green = 8'h53;    Blue = 8'hbe;
end 12'h61a:    begin Red = 8'h07;    Green = 8'h13;    Blue = 8'he4;
end 12'h61b:    begin Red = 8'h6f;    Green = 8'h3e;    Blue = 8'h10;
end 12'h61c:    begin Red = 8'h5b;    Green = 8'h4c;    Blue = 8'h1d;
end 12'h61d:    begin Red = 8'h03;    Green = 8'h42;    Blue = 8'hee;
end 12'h61e:    begin Red = 8'h03;    Green = 8'hf3;    Blue = 8'h7e;
end 12'h61f:    begin Red = 8'hb2;    Green = 8'h7f;    Blue = 8'h48;
end 12'h620:    begin Red = 8'h36;    Green = 8'h34;    Blue = 8'h18;
end 12'h621:    begin Red = 8'hf7;    Green = 8'hbf;    Blue = 8'h9a;
end 12'h622:    begin Red = 8'h3f;    Green = 8'h73;    Blue = 8'h1b;
end 12'h623:    begin Red = 8'hb2;    Green = 8'h63;    Blue = 8'h91;
end 12'h624:    begin Red = 8'hcd;    Green = 8'hce;    Blue = 8'hb9;
end 12'h625:    begin Red = 8'hc5;    Green = 8'he4;    Blue = 8'hd0;
end 12'h626:    begin Red = 8'hce;    Green = 8'h89;    Blue = 8'hb8;
end 12'h627:    begin Red = 8'hc7;    Green = 8'hd5;    Blue = 8'hc6;
end 12'h628:    begin Red = 8'hc4;    Green = 8'hbb;    Blue = 8'h8e;
end 12'h629:    begin Red = 8'h4c;    Green = 8'h68;    Blue = 8'h52;
end 12'h62a:    begin Red = 8'h80;    Green = 8'h7a;    Blue = 8'h16;
end 12'h62b:    begin Red = 8'h08;    Green = 8'h6a;    Blue = 8'h24;
end 12'h62c:    begin Red = 8'h55;    Green = 8'h5e;    Blue = 8'h3b;
end 12'h62d:    begin Red = 8'h07;    Green = 8'he9;    Blue = 8'h6f;
end 12'h62e:    begin Red = 8'h07;    Green = 8'h99;    Blue = 8'h0f;
end 12'h62f:    begin Red = 8'h64;    Green = 8'h83;    Blue = 8'h6b;
end 12'h630:    begin Red = 8'h55;    Green = 8'h81;    Blue = 8'h67;
end 12'h631:    begin Red = 8'h83;    Green = 8'h9b;    Blue = 8'h21;
end 12'h632:    begin Red = 8'h79;    Green = 8'h71;    Blue = 8'h3a;
end 12'h633:    begin Red = 8'hb2;    Green = 8'h73;    Blue = 8'h4c;
end 12'h634:    begin Red = 8'h02;    Green = 8'ha2;    Blue = 8'ha6;
end 12'h635:    begin Red = 8'h03;    Green = 8'hd3;    Blue = 8'h5c;
end 12'h636:    begin Red = 8'h05;    Green = 8'h14;    Blue = 8'hba;
end 12'h637:    begin Red = 8'he9;    Green = 8'hb2;    Blue = 8'h7c;
end 12'h638:    begin Red = 8'he3;    Green = 8'hca;    Blue = 8'h9e;
end 12'h639:    begin Red = 8'h6a;    Green = 8'h50;    Blue = 8'h31;
end 12'h63a:    begin Red = 8'h9e;    Green = 8'h7d;    Blue = 8'h6d;
end 12'h63b:    begin Red = 8'h6b;    Green = 8'h55;    Blue = 8'h1e;
end 12'h63c:    begin Red = 8'h61;    Green = 8'h4b;    Blue = 8'h12;
end 12'h63d:    begin Red = 8'h74;    Green = 8'h4f;    Blue = 8'h36;
end 12'h63e:    begin Red = 8'hcb;    Green = 8'h8a;    Blue = 8'hb3;
end 12'h63f:    begin Red = 8'hc7;    Green = 8'h85;    Blue = 8'hba;
end 12'h640:    begin Red = 8'h85;    Green = 8'ha7;    Blue = 8'h96;
end 12'h641:    begin Red = 8'h5b;    Green = 8'h54;    Blue = 8'h43;
end 12'h642:    begin Red = 8'h66;    Green = 8'h64;    Blue = 8'h37;
end 12'h643:    begin Red = 8'h08;    Green = 8'h49;    Blue = 8'hdf;
end 12'h644:    begin Red = 8'h38;    Green = 8'h4c;    Blue = 8'h11;
end 12'h645:    begin Red = 8'h93;    Green = 8'h61;    Blue = 8'h29;
end 12'h646:    begin Red = 8'h02;    Green = 8'h52;    Blue = 8'h3c;
end 12'h647:    begin Red = 8'h03;    Green = 8'ha3;    Blue = 8'h1d;
end 12'h648:    begin Red = 8'h03;    Green = 8'h52;    Blue = 8'hcd;
end 12'h649:    begin Red = 8'he8;    Green = 8'hb1;    Blue = 8'h82;
end 12'h64a:    begin Red = 8'h72;    Green = 8'h78;    Blue = 8'h4d;
end 12'h64b:    begin Red = 8'h06;    Green = 8'h28;    Blue = 8'h17;
end 12'h64c:    begin Red = 8'h06;    Green = 8'h18;    Blue = 8'h41;
end 12'h64d:    begin Red = 8'h76;    Green = 8'h8f;    Blue = 8'h25;
end 12'h64e:    begin Red = 8'h8f;    Green = 8'h66;    Blue = 8'h2b;
end 12'h64f:    begin Red = 8'h68;    Green = 8'h5b;    Blue = 8'h1e;
end 12'h650:    begin Red = 8'h87;    Green = 8'h59;    Blue = 8'h1e;
end 12'h651:    begin Red = 8'ha7;    Green = 8'ha1;    Blue = 8'h81;
end 12'h652:    begin Red = 8'hc8;    Green = 8'hc0;    Blue = 8'h99;
end 12'h653:    begin Red = 8'ha3;    Green = 8'h9c;    Blue = 8'h83;
end 12'h654:    begin Red = 8'ha1;    Green = 8'h9b;    Blue = 8'h7e;
end 12'h655:    begin Red = 8'hc1;    Green = 8'hb3;    Blue = 8'h20;
end 12'h656:    begin Red = 8'ha8;    Green = 8'hc1;    Blue = 8'h13;
end 12'h657:    begin Red = 8'h13;    Green = 8'h1f;    Blue = 8'h12;
end 12'h658:    begin Red = 8'h68;    Green = 8'h89;    Blue = 8'h12;
end 12'h659:    begin Red = 8'h65;    Green = 8'h90;    Blue = 8'h1a;
end 12'h65a:    begin Red = 8'h8f;    Green = 8'h59;    Blue = 8'h39;
end 12'h65b:    begin Red = 8'h8c;    Green = 8'h58;    Blue = 8'h42;
end 12'h65c:    begin Red = 8'h78;    Green = 8'h96;    Blue = 8'h18;
end 12'h65d:    begin Red = 8'h07;    Green = 8'hd9;    Blue = 8'h2f;
end 12'h65e:    begin Red = 8'h67;    Green = 8'h4c;    Blue = 8'h1b;
end 12'h65f:    begin Red = 8'h59;    Green = 8'h51;    Blue = 8'h1a;
end 12'h660:    begin Red = 8'h6e;    Green = 8'h58;    Blue = 8'h23;
end 12'h661:    begin Red = 8'h77;    Green = 8'h4e;    Blue = 8'h1b;
end 12'h662:    begin Red = 8'hde;    Green = 8'hae;    Blue = 8'h7a;
end 12'h663:    begin Red = 8'h95;    Green = 8'h85;    Blue = 8'h5c;
end 12'h664:    begin Red = 8'h75;    Green = 8'h96;    Blue = 8'h32;
end 12'h665:    begin Red = 8'h05;    Green = 8'hf8;    Blue = 8'h27;
end 12'h666:    begin Red = 8'h05;    Green = 8'hc8;    Blue = 8'h99;
end 12'h667:    begin Red = 8'hff;    Green = 8'he0;    Blue = 8'hbc;
end 12'h668:    begin Red = 8'h66;    Green = 8'h4b;    Blue = 8'h26;
end 12'h669:    begin Red = 8'h03;    Green = 8'h93;    Blue = 8'h5d;
end 12'h66a:    begin Red = 8'h75;    Green = 8'h57;    Blue = 8'h1f;
end 12'h66b:    begin Red = 8'he2;    Green = 8'hd2;    Blue = 8'ha9;
end 12'h66c:    begin Red = 8'had;    Green = 8'ha8;    Blue = 8'h86;
end 12'h66d:    begin Red = 8'ha7;    Green = 8'h96;    Blue = 8'h77;
end 12'h66e:    begin Red = 8'ha8;    Green = 8'hbe;    Blue = 8'h29;
end 12'h66f:    begin Red = 8'h69;    Green = 8'h90;    Blue = 8'h11;
end 12'h670:    begin Red = 8'h71;    Green = 8'h8c;    Blue = 8'h16;
end 12'h671:    begin Red = 8'h72;    Green = 8'h9b;    Blue = 8'h52;
end 12'h672:    begin Red = 8'h55;    Green = 8'h4d;    Blue = 8'h1f;
end 12'h673:    begin Red = 8'h03;    Green = 8'hb3;    Blue = 8'h0e;
end 12'h674:    begin Red = 8'h85;    Green = 8'h78;    Blue = 8'h47;
end 12'h675:    begin Red = 8'h7d;    Green = 8'h8d;    Blue = 8'h1e;
end 12'h676:    begin Red = 8'h70;    Green = 8'h92;    Blue = 8'h15;
end 12'h677:    begin Red = 8'h81;    Green = 8'h71;    Blue = 8'h4e;
end 12'h678:    begin Red = 8'h69;    Green = 8'h50;    Blue = 8'h22;
end 12'h679:    begin Red = 8'h9e;    Green = 8'h6c;    Blue = 8'h33;
end 12'h67a:    begin Red = 8'h85;    Green = 8'h67;    Blue = 8'h2c;
end 12'h67b:    begin Red = 8'h44;    Green = 8'h53;    Blue = 8'h35;
end 12'h67c:    begin Red = 8'h04;    Green = 8'h53;    Blue = 8'h10;
end 12'h67d:    begin Red = 8'hef;    Green = 8'hcd;    Blue = 8'h97;
end 12'h67e:    begin Red = 8'hba;    Green = 8'h62;    Blue = 8'ha1;
end 12'h67f:    begin Red = 8'h60;    Green = 8'h8f;    Blue = 8'h10;
end 12'h680:    begin Red = 8'h88;    Green = 8'h90;    Blue = 8'h20;
end 12'h681:    begin Red = 8'h5b;    Green = 8'h83;    Blue = 8'h46;
end 12'h682:    begin Red = 8'h6a;    Green = 8'ha2;    Blue = 8'h6e;
end 12'h683:    begin Red = 8'h6c;    Green = 8'h98;    Blue = 8'h57;
end 12'h684:    begin Red = 8'h6c;    Green = 8'h99;    Blue = 8'h52;
end 12'h685:    begin Red = 8'h92;    Green = 8'h60;    Blue = 8'h34;
end 12'h686:    begin Red = 8'h52;    Green = 8'h80;    Blue = 8'h48;
end 12'h687:    begin Red = 8'h4e;    Green = 8'h8c;    Blue = 8'h4f;
end 12'h688:    begin Red = 8'h63;    Green = 8'h49;    Blue = 8'h20;
end 12'h689:    begin Red = 8'h04;    Green = 8'h84;    Blue = 8'h5b;
end 12'h68a:    begin Red = 8'hc2;    Green = 8'hb1;    Blue = 8'h8d;
end 12'h68b:    begin Red = 8'h59;    Green = 8'h5d;    Blue = 8'h45;
end 12'h68c:    begin Red = 8'h60;    Green = 8'h65;    Blue = 8'h42;
end 12'h68d:    begin Red = 8'hd5;    Green = 8'hb7;    Blue = 8'h84;
end 12'h68e:    begin Red = 8'hc7;    Green = 8'ha4;    Blue = 8'h77;
end 12'h68f:    begin Red = 8'he4;    Green = 8'hc4;    Blue = 8'h8f;
end 12'h690:    begin Red = 8'hff;    Green = 8'hf3;    Blue = 8'hcc;
end 12'h691:    begin Red = 8'hcc;    Green = 8'hb1;    Blue = 8'h76;
end 12'h692:    begin Red = 8'h97;    Green = 8'h67;    Blue = 8'h23;
end 12'h693:    begin Red = 8'h7e;    Green = 8'h4a;    Blue = 8'h15;
end 12'h694:    begin Red = 8'hae;    Green = 8'hb3;    Blue = 8'h9e;
end 12'h695:    begin Red = 8'h9e;    Green = 8'hb3;    Blue = 8'ha9;
end 12'h696:    begin Red = 8'hbf;    Green = 8'hd4;    Blue = 8'hc9;
end 12'h697:    begin Red = 8'h77;    Green = 8'h6f;    Blue = 8'h5a;
end 12'h698:    begin Red = 8'h7e;    Green = 8'h77;    Blue = 8'h5f;
end 12'h699:    begin Red = 8'h88;    Green = 8'h7f;    Blue = 8'h67;
end 12'h69a:    begin Red = 8'hbd;    Green = 8'hbc;    Blue = 8'h19;
end 12'h69b:    begin Red = 8'h34;    Green = 8'h42;    Blue = 8'h23;
end 12'h69c:    begin Red = 8'h8c;    Green = 8'h8e;    Blue = 8'h2f;
end 12'h69d:    begin Red = 8'hb3;    Green = 8'ha9;    Blue = 8'h2b;
end 12'h69e:    begin Red = 8'hce;    Green = 8'hc7;    Blue = 8'h2d;
end 12'h69f:    begin Red = 8'hc8;    Green = 8'hc2;    Blue = 8'h3c;
end 12'h6a0:    begin Red = 8'h35;    Green = 8'h20;    Blue = 8'h2f;
end 12'h6a1:    begin Red = 8'h09;    Green = 8'h8b;    Blue = 8'h6e;
end 12'h6a2:    begin Red = 8'h8a;    Green = 8'h48;    Blue = 8'h31;
end 12'h6a3:    begin Red = 8'ha6;    Green = 8'h68;    Blue = 8'h2e;
end 12'h6a4:    begin Red = 8'h3a;    Green = 8'h4e;    Blue = 8'h2c;
end 12'h6a5:    begin Red = 8'h06;    Green = 8'hf4;    Blue = 8'h0f;
end 12'h6a6:    begin Red = 8'hd7;    Green = 8'ha7;    Blue = 8'h73;
end 12'h6a7:    begin Red = 8'hb8;    Green = 8'had;    Blue = 8'h83;
end 12'h6a8:    begin Red = 8'hc1;    Green = 8'ha3;    Blue = 8'h6f;
end 12'h6a9:    begin Red = 8'he1;    Green = 8'hc2;    Blue = 8'ha0;
end 12'h6aa:    begin Red = 8'he9;    Green = 8'hcd;    Blue = 8'h97;
end 12'h6ab:    begin Red = 8'h3a;    Green = 8'h4d;    Blue = 8'h31;
end 12'h6ac:    begin Red = 8'he8;    Green = 8'hcf;    Blue = 8'hac;
end 12'h6ad:    begin Red = 8'haf;    Green = 8'h9f;    Blue = 8'ha8;
end 12'h6ae:    begin Red = 8'h6c;    Green = 8'h62;    Blue = 8'h4e;
end 12'h6af:    begin Red = 8'h75;    Green = 8'h6c;    Blue = 8'h53;
end 12'h6b0:    begin Red = 8'hc3;    Green = 8'hab;    Blue = 8'h1a;
end 12'h6b1:    begin Red = 8'h43;    Green = 8'h55;    Blue = 8'h1e;
end 12'h6b2:    begin Red = 8'hc1;    Green = 8'hb5;    Blue = 8'h31;
end 12'h6b3:    begin Red = 8'hba;    Green = 8'ha7;    Blue = 8'h26;
end 12'h6b4:    begin Red = 8'h8d;    Green = 8'had;    Blue = 8'h24;
end 12'h6b5:    begin Red = 8'h72;    Green = 8'h62;    Blue = 8'h21;
end 12'h6b6:    begin Red = 8'h9e;    Green = 8'h65;    Blue = 8'h35;
end 12'h6b7:    begin Red = 8'h53;    Green = 8'h5f;    Blue = 8'h40;
end 12'h6b8:    begin Red = 8'h53;    Green = 8'h5a;    Blue = 8'h41;
end 12'h6b9:    begin Red = 8'h87;    Green = 8'h5c;    Blue = 8'h2a;
end 12'h6ba:    begin Red = 8'h47;    Green = 8'h4d;    Blue = 8'h3c;
end 12'h6bb:    begin Red = 8'h55;    Green = 8'h55;    Blue = 8'h44;
end 12'h6bc:    begin Red = 8'hc8;    Green = 8'ha1;    Blue = 8'h81;
end 12'h6bd:    begin Red = 8'hc4;    Green = 8'hae;    Blue = 8'h88;
end 12'h6be:    begin Red = 8'hb7;    Green = 8'h9f;    Blue = 8'h64;
end 12'h6bf:    begin Red = 8'h72;    Green = 8'h56;    Blue = 8'h13;
end 12'h6c0:    begin Red = 8'h47;    Green = 8'h50;    Blue = 8'h2c;
end 12'h6c1:    begin Red = 8'h4e;    Green = 8'h50;    Blue = 8'h3e;
end 12'h6c2:    begin Red = 8'h81;    Green = 8'h58;    Blue = 8'h25;
end 12'h6c3:    begin Red = 8'hbd;    Green = 8'ha0;    Blue = 8'h69;
end 12'h6c4:    begin Red = 8'hca;    Green = 8'hb8;    Blue = 8'h84;
end 12'h6c5:    begin Red = 8'hcb;    Green = 8'ha8;    Blue = 8'h7d;
end 12'h6c6:    begin Red = 8'hb0;    Green = 8'ha9;    Blue = 8'hab;
end 12'h6c7:    begin Red = 8'h9a;    Green = 8'h91;    Blue = 8'h7c;
end 12'h6c8:    begin Red = 8'h7e;    Green = 8'ha2;    Blue = 8'h6d;
end 12'h6c9:    begin Red = 8'hb8;    Green = 8'ha2;    Blue = 8'h32;
end 12'h6ca:    begin Red = 8'h02;    Green = 8'he2;    Blue = 8'h1e;
end 12'h6cb:    begin Red = 8'h58;    Green = 8'h4d;    Blue = 8'h33;
end 12'h6cc:    begin Red = 8'h05;    Green = 8'ha5;    Blue = 8'h0e;
end 12'h6cd:    begin Red = 8'h9b;    Green = 8'ha2;    Blue = 8'h75;
end 12'h6ce:    begin Red = 8'h26;    Green = 8'h18;    Blue = 8'h17;
end 12'h6cf:    begin Red = 8'h26;    Green = 8'h1b;    Blue = 8'h1e;
end 12'h6d0:    begin Red = 8'h2d;    Green = 8'h1f;    Blue = 8'h1e;
end 12'h6d1:    begin Red = 8'h00;    Green = 8'h10;    Blue = 8'h14;
end 12'h6d2:    begin Red = 8'h31;    Green = 8'h17;    Blue = 8'h1f;
end 12'h6d3:    begin Red = 8'h82;    Green = 8'h9e;    Blue = 8'h68;
end 12'h6d4:    begin Red = 8'h83;    Green = 8'h8c;    Blue = 8'h60;
end 12'h6d5:    begin Red = 8'h7d;    Green = 8'h87;    Blue = 8'h5a;
end 12'h6d6:    begin Red = 8'h7d;    Green = 8'h82;    Blue = 8'h54;
end 12'h6d7:    begin Red = 8'h02;    Green = 8'h4e;    Blue = 8'h1a;
end 12'h6d8:    begin Red = 8'h97;    Green = 8'h8f;    Blue = 8'h75;
end 12'h6d9:    begin Red = 8'h65;    Green = 8'h5d;    Blue = 8'h48;
end 12'h6da:    begin Red = 8'h86;    Green = 8'h9e;    Blue = 8'h77;
end 12'h6db:    begin Red = 8'h35;    Green = 8'h46;    Blue = 8'h14;
end 12'h6dc:    begin Red = 8'h05;    Green = 8'h66;    Blue = 8'h2b;
end 12'h6dd:    begin Red = 8'h63;    Green = 8'h68;    Blue = 8'h1e;
end 12'h6de:    begin Red = 8'h40;    Green = 8'h4a;    Blue = 8'h22;
end 12'h6df:    begin Red = 8'h02;    Green = 8'h23;    Blue = 8'h8b;
end 12'h6e0:    begin Red = 8'hbd;    Green = 8'h7e;    Blue = 8'h49;
end 12'h6e1:    begin Red = 8'h02;    Green = 8'hd2;    Blue = 8'h6a;
end 12'h6e2:    begin Red = 8'h9f;    Green = 8'h68;    Blue = 8'h45;
end 12'h6e3:    begin Red = 8'h00;    Green = 8'h0c;    Blue = 8'h5d;
end 12'h6e4:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h1e;
end 12'h6e5:    begin Red = 8'he9;    Green = 8'hb6;    Blue = 8'h88;
end 12'h6e6:    begin Red = 8'he9;    Green = 8'ha4;    Blue = 8'h77;
end 12'h6e7:    begin Red = 8'h01;    Green = 8'h0b;    Blue = 8'h11;
end 12'h6e8:    begin Red = 8'h83;    Green = 8'h54;    Blue = 8'h16;
end 12'h6e9:    begin Red = 8'haf;    Green = 8'h86;    Blue = 8'h60;
end 12'h6ea:    begin Red = 8'h92;    Green = 8'h99;    Blue = 8'h6a;
end 12'h6eb:    begin Red = 8'h6a;    Green = 8'h6c;    Blue = 8'h4b;
end 12'h6ec:    begin Red = 8'h44;    Green = 8'h31;    Blue = 8'h2c;
end 12'h6ed:    begin Red = 8'he9;    Green = 8'hcc;    Blue = 8'h92;
end 12'h6ee:    begin Red = 8'h4e;    Green = 8'h38;    Blue = 8'h32;
end 12'h6ef:    begin Red = 8'h93;    Green = 8'h9c;    Blue = 8'h61;
end 12'h6f0:    begin Red = 8'h7d;    Green = 8'h53;    Blue = 8'h1d;
end 12'h6f1:    begin Red = 8'hd5;    Green = 8'hbc;    Blue = 8'h87;
end 12'h6f2:    begin Red = 8'hea;    Green = 8'hcb;    Blue = 8'h8c;
end 12'h6f3:    begin Red = 8'h8a;    Green = 8'h82;    Blue = 8'h6f;
end 12'h6f4:    begin Red = 8'h9e;    Green = 8'h96;    Blue = 8'h7e;
end 12'h6f5:    begin Red = 8'h49;    Green = 8'h55;    Blue = 8'h2a;
end 12'h6f6:    begin Red = 8'h03;    Green = 8'h22;    Blue = 8'hdf;
end 12'h6f7:    begin Red = 8'h2b;    Green = 8'h40;    Blue = 8'h12;
end 12'h6f8:    begin Red = 8'h00;    Green = 8'hec;    Blue = 8'h10;
end 12'h6f9:    begin Red = 8'h02;    Green = 8'h21;    Blue = 8'hcf;
end 12'h6fa:    begin Red = 8'h20;    Green = 8'h1b;    Blue = 8'h16;
end 12'h6fb:    begin Red = 8'h85;    Green = 8'h8c;    Blue = 8'h54;
end 12'h6fc:    begin Red = 8'h44;    Green = 8'h48;    Blue = 8'h28;
end 12'h6fd:    begin Red = 8'h73;    Green = 8'h66;    Blue = 8'h54;
end 12'h6fe:    begin Red = 8'ha2;    Green = 8'h85;    Blue = 8'h5e;
end 12'h6ff:    begin Red = 8'haa;    Green = 8'h8e;    Blue = 8'h5c;
end 12'h700:    begin Red = 8'h85;    Green = 8'h77;    Blue = 8'h64;
end 12'h701:    begin Red = 8'h6e;    Green = 8'h5c;    Blue = 8'h50;
end 12'h702:    begin Red = 8'h94;    Green = 8'h86;    Blue = 8'h70;
end 12'h703:    begin Red = 8'h7c;    Green = 8'h6e;    Blue = 8'h64;
end 12'h704:    begin Red = 8'h84;    Green = 8'h92;    Blue = 8'h52;
end 12'h705:    begin Red = 8'h86;    Green = 8'h8c;    Blue = 8'h5a;
end 12'h706:    begin Red = 8'h8e;    Green = 8'h95;    Blue = 8'h5b;
end 12'h707:    begin Red = 8'haf;    Green = 8'h94;    Blue = 8'h5b;
end 12'h708:    begin Red = 8'h86;    Green = 8'h79;    Blue = 8'h5f;
end 12'h709:    begin Red = 8'haf;    Green = 8'hb6;    Blue = 8'hb9;
end 12'h70a:    begin Red = 8'hc5;    Green = 8'hb4;    Blue = 8'h79;
end 12'h70b:    begin Red = 8'hd3;    Green = 8'hc2;    Blue = 8'h84;
end 12'h70c:    begin Red = 8'hb6;    Green = 8'hae;    Blue = 8'h91;
end 12'h70d:    begin Red = 8'hc6;    Green = 8'hbf;    Blue = 8'h9e;
end 12'h70e:    begin Red = 8'h7d;    Green = 8'h9b;    Blue = 8'h74;
end 12'h70f:    begin Red = 8'h03;    Green = 8'hb4;    Blue = 8'h8c;
end 12'h710:    begin Red = 8'h3b;    Green = 8'h46;    Blue = 8'h1e;
end 12'h711:    begin Red = 8'h05;    Green = 8'h96;    Blue = 8'h8f;
end 12'h712:    begin Red = 8'h03;    Green = 8'h72;    Blue = 8'hdd;
end 12'h713:    begin Red = 8'h01;    Green = 8'h62;    Blue = 8'h56;
end 12'h714:    begin Red = 8'hb6;    Green = 8'h7a;    Blue = 8'h4e;
end 12'h715:    begin Red = 8'h02;    Green = 8'ha2;    Blue = 8'h36;
end 12'h716:    begin Red = 8'h75;    Green = 8'h95;    Blue = 8'h78;
end 12'h717:    begin Red = 8'h03;    Green = 8'h14;    Blue = 8'ha4;
end 12'h718:    begin Red = 8'h91;    Green = 8'h6a;    Blue = 8'h3a;
end 12'h719:    begin Red = 8'h59;    Green = 8'h46;    Blue = 8'h31;
end 12'h71a:    begin Red = 8'h99;    Green = 8'ha0;    Blue = 8'h69;
end 12'h71b:    begin Red = 8'h64;    Green = 8'h54;    Blue = 8'h40;
end 12'h71c:    begin Red = 8'h58;    Green = 8'h4d;    Blue = 8'h43;
end 12'h71d:    begin Red = 8'h73;    Green = 8'h66;    Blue = 8'h4c;
end 12'h71e:    begin Red = 8'h84;    Green = 8'h8f;    Blue = 8'h48;
end 12'h71f:    begin Red = 8'hee;    Green = 8'hd9;    Blue = 8'had;
end 12'h720:    begin Red = 8'h83;    Green = 8'h73;    Blue = 8'h54;
end 12'h721:    begin Red = 8'h78;    Green = 8'h69;    Blue = 8'h5a;
end 12'h722:    begin Red = 8'hc9;    Green = 8'hc7;    Blue = 8'hca;
end 12'h723:    begin Red = 8'hca;    Green = 8'hb9;    Blue = 8'h7e;
end 12'h724:    begin Red = 8'hbc;    Green = 8'haf;    Blue = 8'h77;
end 12'h725:    begin Red = 8'had;    Green = 8'ha7;    Blue = 8'h8b;
end 12'h726:    begin Red = 8'hb5;    Green = 8'hac;    Blue = 8'h8c;
end 12'h727:    begin Red = 8'h8e;    Green = 8'hb2;    Blue = 8'h8a;
end 12'h728:    begin Red = 8'h51;    Green = 8'h61;    Blue = 8'h2a;
end 12'h729:    begin Red = 8'h48;    Green = 8'h5f;    Blue = 8'h2b;
end 12'h72a:    begin Red = 8'h04;    Green = 8'h63;    Blue = 8'h8e;
end 12'h72b:    begin Red = 8'h77;    Green = 8'h65;    Blue = 8'h36;
end 12'h72c:    begin Red = 8'h02;    Green = 8'h62;    Blue = 8'hd9;
end 12'h72d:    begin Red = 8'h6b;    Green = 8'h8e;    Blue = 8'h7a;
end 12'h72e:    begin Red = 8'h04;    Green = 8'h55;    Blue = 8'h4e;
end 12'h72f:    begin Red = 8'h97;    Green = 8'h68;    Blue = 8'h36;
end 12'h730:    begin Red = 8'h63;    Green = 8'h39;    Blue = 8'h23;
end 12'h731:    begin Red = 8'h92;    Green = 8'h9a;    Blue = 8'h5c;
end 12'h732:    begin Red = 8'hd8;    Green = 8'hcf;    Blue = 8'h96;
end 12'h733:    begin Red = 8'h5e;    Green = 8'h4f;    Blue = 8'h43;
end 12'h734:    begin Red = 8'h44;    Green = 8'h52;    Blue = 8'h76;
end 12'h735:    begin Red = 8'h3f;    Green = 8'h54;    Blue = 8'h81;
end 12'h736:    begin Red = 8'h47;    Green = 8'h58;    Blue = 8'h7b;
end 12'h737:    begin Red = 8'h70;    Green = 8'h99;    Blue = 8'he2;
end 12'h738:    begin Red = 8'h65;    Green = 8'h58;    Blue = 8'h48;
end 12'h739:    begin Red = 8'h66;    Green = 8'h58;    Blue = 8'h4d;
end 12'h73a:    begin Red = 8'h4b;    Green = 8'h66;    Blue = 8'h91;
end 12'h73b:    begin Red = 8'h4f;    Green = 8'h5f;    Blue = 8'h91;
end 12'h73c:    begin Red = 8'h91;    Green = 8'ha7;    Blue = 8'he7;
end 12'h73d:    begin Red = 8'h7f;    Green = 8'ha4;    Blue = 8'hed;
end 12'h73e:    begin Red = 8'h49;    Green = 8'h5e;    Blue = 8'h89;
end 12'h73f:    begin Red = 8'h50;    Green = 8'h62;    Blue = 8'h86;
end 12'h740:    begin Red = 8'h90;    Green = 8'h95;    Blue = 8'h47;
end 12'h741:    begin Red = 8'he6;    Green = 8'hc0;    Blue = 8'h89;
end 12'h742:    begin Red = 8'h3e;    Green = 8'h52;    Blue = 8'h7a;
end 12'h743:    begin Red = 8'h41;    Green = 8'h56;    Blue = 8'h8b;
end 12'h744:    begin Red = 8'h71;    Green = 8'h8d;    Blue = 8'hd0;
end 12'h745:    begin Red = 8'hbd;    Green = 8'h75;    Blue = 8'haa;
end 12'h746:    begin Red = 8'hb8;    Green = 8'h64;    Blue = 8'h96;
end 12'h747:    begin Red = 8'h84;    Green = 8'h74;    Blue = 8'h6a;
end 12'h748:    begin Red = 8'hdd;    Green = 8'hcc;    Blue = 8'ha7;
end 12'h749:    begin Red = 8'h8b;    Green = 8'h7c;    Blue = 8'h70;
end 12'h74a:    begin Red = 8'hcf;    Green = 8'hbd;    Blue = 8'h7f;
end 12'h74b:    begin Red = 8'h04;    Green = 8'h13;    Blue = 8'h4e;
end 12'h74c:    begin Red = 8'h45;    Green = 8'h2f;    Blue = 8'h1a;
end 12'h74d:    begin Red = 8'h03;    Green = 8'h32;    Blue = 8'ha9;
end 12'h74e:    begin Red = 8'h00;    Green = 8'h13;    Blue = 8'hff;
end 12'h74f:    begin Red = 8'h1d;    Green = 8'h1a;    Blue = 8'h10;
end 12'h750:    begin Red = 8'h2f;    Green = 8'h25;    Blue = 8'h1a;
end 12'h751:    begin Red = 8'h73;    Green = 8'h61;    Blue = 8'h44;
end 12'h752:    begin Red = 8'hd3;    Green = 8'ha5;    Blue = 8'h7c;
end 12'h753:    begin Red = 8'hc6;    Green = 8'h8e;    Blue = 8'h5e;
end 12'h754:    begin Red = 8'h69;    Green = 8'h6f;    Blue = 8'h42;
end 12'h755:    begin Red = 8'he3;    Green = 8'hd9;    Blue = 8'ha4;
end 12'h756:    begin Red = 8'hd3;    Green = 8'hd8;    Blue = 8'haa;
end 12'h757:    begin Red = 8'h50;    Green = 8'h53;    Blue = 8'h39;
end 12'h758:    begin Red = 8'hea;    Green = 8'he1;    Blue = 8'hb1;
end 12'h759:    begin Red = 8'haf;    Green = 8'ha7;    Blue = 8'h75;
end 12'h75a:    begin Red = 8'hae;    Green = 8'ha4;    Blue = 8'h7e;
end 12'h75b:    begin Red = 8'h60;    Green = 8'h58;    Blue = 8'h47;
end 12'h75c:    begin Red = 8'h8b;    Green = 8'h6b;    Blue = 8'h4d;
end 12'h75d:    begin Red = 8'h83;    Green = 8'h97;    Blue = 8'h55;
end 12'h75e:    begin Red = 8'h65;    Green = 8'h53;    Blue = 8'h49;
end 12'h75f:    begin Red = 8'hb7;    Green = 8'h73;    Blue = 8'hb1;
end 12'h760:    begin Red = 8'hdb;    Green = 8'h86;    Blue = 8'hbe;
end 12'h761:    begin Red = 8'hc9;    Green = 8'h81;    Blue = 8'hbf;
end 12'h762:    begin Red = 8'hd2;    Green = 8'h7f;    Blue = 8'hba;
end 12'h763:    begin Red = 8'hb3;    Green = 8'ha6;    Blue = 8'h6c;
end 12'h764:    begin Red = 8'hb9;    Green = 8'had;    Blue = 8'h70;
end 12'h765:    begin Red = 8'haf;    Green = 8'ha1;    Blue = 8'h77;
end 12'h766:    begin Red = 8'h87;    Green = 8'h73;    Blue = 8'h76;
end 12'h767:    begin Red = 8'h7c;    Green = 8'h67;    Blue = 8'h65;
end 12'h768:    begin Red = 8'hcd;    Green = 8'hc0;    Blue = 8'h85;
end 12'h769:    begin Red = 8'h8c;    Green = 8'hb1;    Blue = 8'h99;
end 12'h76a:    begin Red = 8'h36;    Green = 8'h47;    Blue = 8'h21;
end 12'h76b:    begin Red = 8'h02;    Green = 8'he2;    Blue = 8'ha4;
end 12'h76c:    begin Red = 8'h6b;    Green = 8'h62;    Blue = 8'h21;
end 12'h76d:    begin Red = 8'h37;    Green = 8'h2a;    Blue = 8'h16;
end 12'h76e:    begin Red = 8'h73;    Green = 8'h6c;    Blue = 8'h39;
end 12'h76f:    begin Red = 8'h03;    Green = 8'h73;    Blue = 8'h1c;
end 12'h770:    begin Red = 8'h71;    Green = 8'h51;    Blue = 8'h23;
end 12'h771:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h9e;
end 12'h772:    begin Red = 8'h02;    Green = 8'hd2;    Blue = 8'h9e;
end 12'h773:    begin Red = 8'h5c;    Green = 8'h4a;    Blue = 8'h12;
end 12'h774:    begin Red = 8'ha5;    Green = 8'h78;    Blue = 8'h4f;
end 12'h775:    begin Red = 8'h7e;    Green = 8'h5a;    Blue = 8'h31;
end 12'h776:    begin Red = 8'h00;    Green = 8'h12;    Blue = 8'hee;
end 12'h777:    begin Red = 8'hdb;    Green = 8'had;    Blue = 8'h83;
end 12'h778:    begin Red = 8'hdd;    Green = 8'ha3;    Blue = 8'h70;
end 12'h779:    begin Red = 8'hc3;    Green = 8'hb9;    Blue = 8'h88;
end 12'h77a:    begin Red = 8'ha8;    Green = 8'h9e;    Blue = 8'h78;
end 12'h77b:    begin Red = 8'h7f;    Green = 8'h68;    Blue = 8'h58;
end 12'h77c:    begin Red = 8'h7e;    Green = 8'h6b;    Blue = 8'h5f;
end 12'h77d:    begin Red = 8'h6e;    Green = 8'h5a;    Blue = 8'h49;
end 12'h77e:    begin Red = 8'h85;    Green = 8'h7a;    Blue = 8'h6d;
end 12'h77f:    begin Red = 8'h90;    Green = 8'h72;    Blue = 8'h62;
end 12'h780:    begin Red = 8'h75;    Green = 8'h66;    Blue = 8'h63;
end 12'h781:    begin Red = 8'h5a;    Green = 8'h5c;    Blue = 8'h3e;
end 12'h782:    begin Red = 8'hd3;    Green = 8'h8e;    Blue = 8'hbe;
end 12'h783:    begin Red = 8'hb0;    Green = 8'ha1;    Blue = 8'h72;
end 12'h784:    begin Red = 8'ha8;    Green = 8'h9a;    Blue = 8'h6e;
end 12'h785:    begin Red = 8'h82;    Green = 8'h6f;    Blue = 8'h6a;
end 12'h786:    begin Red = 8'h41;    Green = 8'h42;    Blue = 8'h11;
end 12'h787:    begin Red = 8'h79;    Green = 8'h90;    Blue = 8'h2b;
end 12'h788:    begin Red = 8'h96;    Green = 8'h5b;    Blue = 8'h2b;
end 12'h789:    begin Red = 8'haa;    Green = 8'h78;    Blue = 8'h4d;
end 12'h78a:    begin Red = 8'h03;    Green = 8'he3;    Blue = 8'h25;
end 12'h78b:    begin Red = 8'h05;    Green = 8'h24;    Blue = 8'h9c;
end 12'h78c:    begin Red = 8'h97;    Green = 8'h65;    Blue = 8'h3c;
end 12'h78d:    begin Red = 8'h3d;    Green = 8'h59;    Blue = 8'h74;
end 12'h78e:    begin Red = 8'h43;    Green = 8'h59;    Blue = 8'h81;
end 12'h78f:    begin Red = 8'h7e;    Green = 8'ha2;    Blue = 8'he7;
end 12'h790:    begin Red = 8'h76;    Green = 8'h90;    Blue = 8'hd5;
end 12'h791:    begin Red = 8'h4e;    Green = 8'h62;    Blue = 8'h8b;
end 12'h792:    begin Red = 8'h4d;    Green = 8'h61;    Blue = 8'h9c;
end 12'h793:    begin Red = 8'h85;    Green = 8'ha7;    Blue = 8'heb;
end 12'h794:    begin Red = 8'h7b;    Green = 8'ha8;    Blue = 8'he8;
end 12'h795:    begin Red = 8'h82;    Green = 8'had;    Blue = 8'hea;
end 12'h796:    begin Red = 8'h7b;    Green = 8'h6b;    Blue = 8'h43;
end 12'h797:    begin Red = 8'h86;    Green = 8'ha7;    Blue = 8'hf2;
end 12'h798:    begin Red = 8'h93;    Green = 8'hb8;    Blue = 8'hf4;
end 12'h799:    begin Red = 8'h4e;    Green = 8'h64;    Blue = 8'h96;
end 12'h79a:    begin Red = 8'h55;    Green = 8'h62;    Blue = 8'h8f;
end 12'h79b:    begin Red = 8'h78;    Green = 8'h9d;    Blue = 8'he2;
end 12'h79c:    begin Red = 8'hd8;    Green = 8'hc8;    Blue = 8'haa;
end 12'h79d:    begin Red = 8'he1;    Green = 8'hd1;    Blue = 8'hb2;
end 12'h79e:    begin Red = 8'h02;    Green = 8'h22;    Blue = 8'h97;
end 12'h79f:    begin Red = 8'h8c;    Green = 8'ha5;    Blue = 8'h23;
end 12'h7a0:    begin Red = 8'h8e;    Green = 8'h68;    Blue = 8'h24;
end 12'h7a1:    begin Red = 8'h5d;    Green = 8'h6e;    Blue = 8'h45;
end 12'h7a2:    begin Red = 8'h77;    Green = 8'h7e;    Blue = 8'h4d;
end 12'h7a3:    begin Red = 8'hdf;    Green = 8'hd7;    Blue = 8'h98;
end 12'h7a4:    begin Red = 8'he8;    Green = 8'hde;    Blue = 8'hac;
end 12'h7a5:    begin Red = 8'h39;    Green = 8'h59;    Blue = 8'h79;
end 12'h7a6:    begin Red = 8'h47;    Green = 8'h56;    Blue = 8'h8d;
end 12'h7a7:    begin Red = 8'h79;    Green = 8'h9f;    Blue = 8'hee;
end 12'h7a8:    begin Red = 8'h6f;    Green = 8'h91;    Blue = 8'he3;
end 12'h7a9:    begin Red = 8'h79;    Green = 8'h92;    Blue = 8'hd0;
end 12'h7aa:    begin Red = 8'h87;    Green = 8'h6a;    Blue = 8'h42;
end 12'h7ab:    begin Red = 8'h65;    Green = 8'h69;    Blue = 8'h48;
end 12'h7ac:    begin Red = 8'h6f;    Green = 8'h94;    Blue = 8'hd9;
end 12'h7ad:    begin Red = 8'h6a;    Green = 8'h93;    Blue = 8'hd3;
end 12'h7ae:    begin Red = 8'ha2;    Green = 8'had;    Blue = 8'h9f;
end 12'h7af:    begin Red = 8'h7b;    Green = 8'h6a;    Blue = 8'h6a;
end 12'h7b0:    begin Red = 8'h07;    Green = 8'h68;    Blue = 8'hfe;
end 12'h7b1:    begin Red = 8'h01;    Green = 8'hb1;    Blue = 8'hcc;
end 12'h7b2:    begin Red = 8'h00;    Green = 8'h09;    Blue = 8'h86;
end 12'h7b3:    begin Red = 8'h00;    Green = 8'hf1;    Blue = 8'h35;
end 12'h7b4:    begin Red = 8'h8a;    Green = 8'ha4;    Blue = 8'h2a;
end 12'h7b5:    begin Red = 8'h99;    Green = 8'hb5;    Blue = 8'h33;
end 12'h7b6:    begin Red = 8'h73;    Green = 8'h5c;    Blue = 8'h22;
end 12'h7b7:    begin Red = 8'h03;    Green = 8'h62;    Blue = 8'h65;
end 12'h7b8:    begin Red = 8'h02;    Green = 8'hd2;    Blue = 8'h1b;
end 12'h7b9:    begin Red = 8'h84;    Green = 8'h4f;    Blue = 8'h16;
end 12'h7ba:    begin Red = 8'h07;    Green = 8'hc4;    Blue = 8'h4e;
end 12'h7bb:    begin Red = 8'h70;    Green = 8'h86;    Blue = 8'h50;
end 12'h7bc:    begin Red = 8'h9b;    Green = 8'h94;    Blue = 8'h72;
end 12'h7bd:    begin Red = 8'hc8;    Green = 8'hcc;    Blue = 8'h9b;
end 12'h7be:    begin Red = 8'h92;    Green = 8'h92;    Blue = 8'h6b;
end 12'h7bf:    begin Red = 8'h79;    Green = 8'h71;    Blue = 8'h53;
end 12'h7c0:    begin Red = 8'h50;    Green = 8'h65;    Blue = 8'h90;
end 12'h7c1:    begin Red = 8'h5e;    Green = 8'h53;    Blue = 8'h48;
end 12'h7c2:    begin Red = 8'hac;    Green = 8'hb4;    Blue = 8'h99;
end 12'h7c3:    begin Red = 8'hcd;    Green = 8'h90;    Blue = 8'hba;
end 12'h7c4:    begin Red = 8'h31;    Green = 8'h30;    Blue = 8'h16;
end 12'h7c5:    begin Red = 8'h02;    Green = 8'h32;    Blue = 8'h8a;
end 12'h7c6:    begin Red = 8'h45;    Green = 8'h4b;    Blue = 8'h18;
end 12'h7c7:    begin Red = 8'h8d;    Green = 8'h61;    Blue = 8'h2d;
end 12'h7c8:    begin Red = 8'h98;    Green = 8'h7f;    Blue = 8'h4f;
end 12'h7c9:    begin Red = 8'h01;    Green = 8'h1f;    Blue = 8'h13;
end 12'h7ca:    begin Red = 8'h01;    Green = 8'ha1;    Blue = 8'h8c;
end 12'h7cb:    begin Red = 8'h31;    Green = 8'h2a;    Blue = 8'h17;
end 12'h7cc:    begin Red = 8'h57;    Green = 8'h6d;    Blue = 8'h42;
end 12'h7cd:    begin Red = 8'h2f;    Green = 8'h24;    Blue = 8'h1f;
end 12'h7ce:    begin Red = 8'hac;    Green = 8'hb3;    Blue = 8'h83;
end 12'h7cf:    begin Red = 8'h97;    Green = 8'h9e;    Blue = 8'h6f;
end 12'h7d0:    begin Red = 8'hbe;    Green = 8'h71;    Blue = 8'h9b;
end 12'h7d1:    begin Red = 8'hab;    Green = 8'h64;    Blue = 8'h9e;
end 12'h7d2:    begin Red = 8'hc8;    Green = 8'hbc;    Blue = 8'hc2;
end 12'h7d3:    begin Red = 8'h87;    Green = 8'h74;    Blue = 8'h6f;
end 12'h7d4:    begin Red = 8'hd6;    Green = 8'hc7;    Blue = 8'h97;
end 12'h7d5:    begin Red = 8'hb7;    Green = 8'ha2;    Blue = 8'h8e;
end 12'h7d6:    begin Red = 8'h81;    Green = 8'hb4;    Blue = 8'h93;
end 12'h7d7:    begin Red = 8'h6c;    Green = 8'h69;    Blue = 8'h1c;
end 12'h7d8:    begin Red = 8'h62;    Green = 8'h5f;    Blue = 8'h14;
end 12'h7d9:    begin Red = 8'h7b;    Green = 8'h98;    Blue = 8'h48;
end 12'h7da:    begin Red = 8'h6d;    Green = 8'h88;    Blue = 8'h34;
end 12'h7db:    begin Red = 8'h31;    Green = 8'h2e;    Blue = 8'h21;
end 12'h7dc:    begin Red = 8'h3d;    Green = 8'h53;    Blue = 8'h1d;
end 12'h7dd:    begin Red = 8'h06;    Green = 8'h14;    Blue = 8'h76;
end 12'h7de:    begin Red = 8'h77;    Green = 8'h46;    Blue = 8'h16;
end 12'h7df:    begin Red = 8'h72;    Green = 8'h74;    Blue = 8'h55;
end 12'h7e0:    begin Red = 8'h83;    Green = 8'h83;    Blue = 8'h61;
end 12'h7e1:    begin Red = 8'hb9;    Green = 8'h74;    Blue = 8'ha2;
end 12'h7e2:    begin Red = 8'hc1;    Green = 8'hc6;    Blue = 8'hc9;
end 12'h7e3:    begin Red = 8'hb1;    Green = 8'hac;    Blue = 8'h73;
end 12'h7e4:    begin Red = 8'hb7;    Green = 8'haf;    Blue = 8'h7d;
end 12'h7e5:    begin Red = 8'hd8;    Green = 8'hc4;    Blue = 8'h8f;
end 12'h7e6:    begin Red = 8'h58;    Green = 8'h4e;    Blue = 8'h2c;
end 12'h7e7:    begin Red = 8'h6f;    Green = 8'h88;    Blue = 8'h3b;
end 12'h7e8:    begin Red = 8'h2c;    Green = 8'h2f;    Blue = 8'h1e;
end 12'h7e9:    begin Red = 8'ha1;    Green = 8'h63;    Blue = 8'h2a;
end 12'h7ea:    begin Red = 8'h7e;    Green = 8'h5a;    Blue = 8'h1a;
end 12'h7eb:    begin Red = 8'h9e;    Green = 8'h75;    Blue = 8'h59;
end 12'h7ec:    begin Red = 8'h83;    Green = 8'h98;    Blue = 8'h6c;
end 12'h7ed:    begin Red = 8'h6c;    Green = 8'h65;    Blue = 8'h17;
end 12'h7ee:    begin Red = 8'h4c;    Green = 8'h4a;    Blue = 8'h1e;
end 12'h7ef:    begin Red = 8'h7f;    Green = 8'h52;    Blue = 8'h2c;
end 12'h7f0:    begin Red = 8'h05;    Green = 8'h84;    Blue = 8'hd6;
end 12'h7f1:    begin Red = 8'h06;    Green = 8'h05;    Blue = 8'h5e;
end 12'h7f2:    begin Red = 8'h90;    Green = 8'h5e;    Blue = 8'h3c;
end 12'h7f3:    begin Red = 8'hc1;    Green = 8'h93;    Blue = 8'h61;
end 12'h7f4:    begin Red = 8'hbe;    Green = 8'h8c;    Blue = 8'h64;
end 12'h7f5:    begin Red = 8'hae;    Green = 8'h64;    Blue = 8'h97;
end 12'h7f6:    begin Red = 8'hca;    Green = 8'hde;    Blue = 8'hcc;
end 12'h7f7:    begin Red = 8'hc8;    Green = 8'h84;    Blue = 8'hb5;
end 12'h7f8:    begin Red = 8'h8a;    Green = 8'h7c;    Blue = 8'h1c;
end 12'h7f9:    begin Red = 8'h73;    Green = 8'h6b;    Blue = 8'h1d;
end 12'h7fa:    begin Red = 8'h61;    Green = 8'h6a;    Blue = 8'h14;
end 12'h7fb:    begin Red = 8'h69;    Green = 8'h88;    Blue = 8'h18;
end 12'h7fc:    begin Red = 8'h03;    Green = 8'h64;    Blue = 8'hf6;
end 12'h7fd:    begin Red = 8'h83;    Green = 8'h91;    Blue = 8'h63;
end 12'h7fe:    begin Red = 8'h89;    Green = 8'h4c;    Blue = 8'h1a;
end 12'h7ff:    begin Red = 8'h5b;    Green = 8'h87;    Blue = 8'h68;
end 12'h800:    begin Red = 8'h5e;    Green = 8'h88;    Blue = 8'h77;
end 12'h801:    begin Red = 8'h79;    Green = 8'h53;    Blue = 8'h26;
end 12'h802:    begin Red = 8'h61;    Green = 8'h88;    Blue = 8'h80;
end 12'h803:    begin Red = 8'h9d;    Green = 8'h81;    Blue = 8'h4a;
end 12'h804:    begin Red = 8'ha0;    Green = 8'ha6;    Blue = 8'h75;
end 12'h805:    begin Red = 8'hc9;    Green = 8'hcc;    Blue = 8'ha0;
end 12'h806:    begin Red = 8'hb2;    Green = 8'h5c;    Blue = 8'h99;
end 12'h807:    begin Red = 8'h77;    Green = 8'h7c;    Blue = 8'h1c;
end 12'h808:    begin Red = 8'h72;    Green = 8'h6b;    Blue = 8'h13;
end 12'h809:    begin Red = 8'h05;    Green = 8'hc6;    Blue = 8'haf;
end 12'h80a:    begin Red = 8'h63;    Green = 8'h7e;    Blue = 8'h17;
end 12'h80b:    begin Red = 8'h04;    Green = 8'h04;    Blue = 8'hfe;
end 12'h80c:    begin Red = 8'h03;    Green = 8'h94;    Blue = 8'hd9;
end 12'h80d:    begin Red = 8'h5a;    Green = 8'h82;    Blue = 8'h6d;
end 12'h80e:    begin Red = 8'ha5;    Green = 8'h8a;    Blue = 8'h53;
end 12'h80f:    begin Red = 8'ha5;    Green = 8'h78;    Blue = 8'h5b;
end 12'h810:    begin Red = 8'hac;    Green = 8'hb0;    Blue = 8'h89;
end 12'h811:    begin Red = 8'h7e;    Green = 8'h78;    Blue = 8'h59;
end 12'h812:    begin Red = 8'h8b;    Green = 8'ha8;    Blue = 8'h95;
end 12'h813:    begin Red = 8'h7e;    Green = 8'h6c;    Blue = 8'h10;
end 12'h814:    begin Red = 8'h77;    Green = 8'h70;    Blue = 8'h1c;
end 12'h815:    begin Red = 8'h51;    Green = 8'h4d;    Blue = 8'h18;
end 12'h816:    begin Red = 8'h04;    Green = 8'hd6;    Blue = 8'h39;
end 12'h817:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'hbc;
end 12'h818:    begin Red = 8'h00;    Green = 8'h08;    Blue = 8'ha7;
end 12'h819:    begin Red = 8'ha2;    Green = 8'h5e;    Blue = 8'h33;
end 12'h81a:    begin Red = 8'h4b;    Green = 8'h7d;    Blue = 8'h44;
end 12'h81b:    begin Red = 8'h5c;    Green = 8'h92;    Blue = 8'h52;
end 12'h81c:    begin Red = 8'h5f;    Green = 8'h8d;    Blue = 8'h50;
end 12'h81d:    begin Red = 8'h5f;    Green = 8'h8c;    Blue = 8'h44;
end 12'h81e:    begin Red = 8'hc8;    Green = 8'hd6;    Blue = 8'hab;
end 12'h81f:    begin Red = 8'hdc;    Green = 8'he1;    Blue = 8'hb1;
end 12'h820:    begin Red = 8'h46;    Green = 8'h7f;    Blue = 8'h43;
end 12'h821:    begin Red = 8'h48;    Green = 8'h76;    Blue = 8'h3e;
end 12'h822:    begin Red = 8'h88;    Green = 8'h8a;    Blue = 8'h67;
end 12'h823:    begin Red = 8'h74;    Green = 8'h91;    Blue = 8'hdb;
end 12'h824:    begin Red = 8'hcd;    Green = 8'hd2;    Blue = 8'ha4;
end 12'h825:    begin Red = 8'hb3;    Green = 8'h45;    Blue = 8'h90;
end 12'h826:    begin Red = 8'hcc;    Green = 8'hd9;    Blue = 8'hd1;
end 12'h827:    begin Red = 8'hac;    Green = 8'ha3;    Blue = 8'h86;
end 12'h828:    begin Red = 8'h06;    Green = 8'hd5;    Blue = 8'hf0;
end 12'h829:    begin Red = 8'h06;    Green = 8'h36;    Blue = 8'h6f;
end 12'h82a:    begin Red = 8'h06;    Green = 8'ha8;    Blue = 8'he5;
end 12'h82b:    begin Red = 8'h03;    Green = 8'ha4;    Blue = 8'h9c;
end 12'h82c:    begin Red = 8'h69;    Green = 8'h83;    Blue = 8'h10;
end 12'h82d:    begin Red = 8'h00;    Green = 8'h15;    Blue = 8'he8;
end 12'h82e:    begin Red = 8'h05;    Green = 8'h87;    Blue = 8'h4b;
end 12'h82f:    begin Red = 8'h00;    Green = 8'h0a;    Blue = 8'hd4;
end 12'h830:    begin Red = 8'h67;    Green = 8'h98;    Blue = 8'h52;
end 12'h831:    begin Red = 8'h61;    Green = 8'h94;    Blue = 8'h4d;
end 12'h832:    begin Red = 8'h67;    Green = 8'h92;    Blue = 8'h58;
end 12'h833:    begin Red = 8'he2;    Green = 8'he7;    Blue = 8'hbc;
end 12'h834:    begin Red = 8'hb4;    Green = 8'ha6;    Blue = 8'ha6;
end 12'h835:    begin Red = 8'h05;    Green = 8'h66;    Blue = 8'h3e;
end 12'h836:    begin Red = 8'h53;    Green = 8'h5e;    Blue = 8'h12;
end 12'h837:    begin Red = 8'h3f;    Green = 8'h40;    Blue = 8'h19;
end 12'h838:    begin Red = 8'h60;    Green = 8'h78;    Blue = 8'h10;
end 12'h839:    begin Red = 8'h66;    Green = 8'h7c;    Blue = 8'h10;
end 12'h83a:    begin Red = 8'h01;    Green = 8'h21;    Blue = 8'h26;
end 12'h83b:    begin Red = 8'h01;    Green = 8'hb2;    Blue = 8'h5a;
end 12'h83c:    begin Red = 8'h01;    Green = 8'h51;    Blue = 8'he0;
end 12'h83d:    begin Red = 8'h9d;    Green = 8'h5e;    Blue = 8'h38;
end 12'h83e:    begin Red = 8'h55;    Green = 8'h7a;    Blue = 8'h46;
end 12'h83f:    begin Red = 8'ha5;    Green = 8'hba;    Blue = 8'h8d;
end 12'h840:    begin Red = 8'h7e;    Green = 8'h73;    Blue = 8'h3f;
end 12'h841:    begin Red = 8'h95;    Green = 8'h99;    Blue = 8'h73;
end 12'h842:    begin Red = 8'hee;    Green = 8'hd3;    Blue = 8'h98;
end 12'h843:    begin Red = 8'hae;    Green = 8'h51;    Blue = 8'h9a;
end 12'h844:    begin Red = 8'h54;    Green = 8'h43;    Blue = 8'h2b;
end 12'h845:    begin Red = 8'h63;    Green = 8'h41;    Blue = 8'h2d;
end 12'h846:    begin Red = 8'h6d;    Green = 8'h42;    Blue = 8'h31;
end 12'h847:    begin Red = 8'h86;    Green = 8'hb1;    Blue = 8'hb0;
end 12'h848:    begin Red = 8'h8f;    Green = 8'h87;    Blue = 8'h13;
end 12'h849:    begin Red = 8'h72;    Green = 8'h71;    Blue = 8'h17;
end 12'h84a:    begin Red = 8'h22;    Green = 8'h10;    Blue = 8'h1d;
end 12'h84b:    begin Red = 8'h02;    Green = 8'h0f;    Blue = 8'h20;
end 12'h84c:    begin Red = 8'h40;    Green = 8'h1c;    Blue = 8'h1d;
end 12'h84d:    begin Red = 8'h05;    Green = 8'h06;    Blue = 8'h1f;
end 12'h84e:    begin Red = 8'h3f;    Green = 8'h29;    Blue = 8'h1d;
end 12'h84f:    begin Red = 8'h02;    Green = 8'he2;    Blue = 8'hed;
end 12'h850:    begin Red = 8'h02;    Green = 8'h52;    Blue = 8'hff;
end 12'h851:    begin Red = 8'h01;    Green = 8'h21;    Blue = 8'h71;
end 12'h852:    begin Red = 8'h93;    Green = 8'hb3;    Blue = 8'h8f;
end 12'h853:    begin Red = 8'h5e;    Green = 8'h87;    Blue = 8'h51;
end 12'h854:    begin Red = 8'h76;    Green = 8'ha7;    Blue = 8'h64;
end 12'h855:    begin Red = 8'h70;    Green = 8'ha0;    Blue = 8'h62;
end 12'h856:    begin Red = 8'h59;    Green = 8'h84;    Blue = 8'h4d;
end 12'h857:    begin Red = 8'h85;    Green = 8'h7a;    Blue = 8'h55;
end 12'h858:    begin Red = 8'h76;    Green = 8'h60;    Blue = 8'h59;
end 12'h859:    begin Red = 8'hca;    Green = 8'hcc;    Blue = 8'hd0;
end 12'h85a:    begin Red = 8'h07;    Green = 8'h86;    Blue = 8'h79;
end 12'h85b:    begin Red = 8'h86;    Green = 8'h86;    Blue = 8'h20;
end 12'h85c:    begin Red = 8'h78;    Green = 8'h76;    Blue = 8'h1c;
end 12'h85d:    begin Red = 8'h27;    Green = 8'h21;    Blue = 8'h14;
end 12'h85e:    begin Red = 8'h01;    Green = 8'hb1;    Blue = 8'h7e;
end 12'h85f:    begin Red = 8'h4f;    Green = 8'h63;    Blue = 8'h16;
end 12'h860:    begin Red = 8'h02;    Green = 8'h53;    Blue = 8'h09;
end 12'h861:    begin Red = 8'h97;    Green = 8'h5c;    Blue = 8'h36;
end 12'h862:    begin Red = 8'hcb;    Green = 8'hdb;    Blue = 8'hb1;
end 12'h863:    begin Red = 8'h7d;    Green = 8'h60;    Blue = 8'h5d;
end 12'h864:    begin Red = 8'h02;    Green = 8'hc3;    Blue = 8'h99;
end 12'h865:    begin Red = 8'ha3;    Green = 8'hb3;    Blue = 8'h8a;
end 12'h866:    begin Red = 8'hb9;    Green = 8'hbe;    Blue = 8'h92;
end 12'h867:    begin Red = 8'ha9;    Green = 8'hae;    Blue = 8'h80;
end 12'h868:    begin Red = 8'h32;    Green = 8'h53;    Blue = 8'h80;
end 12'h869:    begin Red = 8'h35;    Green = 8'h50;    Blue = 8'h8b;
end 12'h86a:    begin Red = 8'h2f;    Green = 8'h50;    Blue = 8'h8b;
end 12'h86b:    begin Red = 8'h3a;    Green = 8'h4f;    Blue = 8'h87;
end 12'h86c:    begin Red = 8'h6c;    Green = 8'h56;    Blue = 8'h4f;
end 12'h86d:    begin Red = 8'h3d;    Green = 8'h5c;    Blue = 8'h8b;
end 12'h86e:    begin Red = 8'h44;    Green = 8'h5c;    Blue = 8'h9b;
end 12'h86f:    begin Red = 8'h3e;    Green = 8'h5b;    Blue = 8'h9d;
end 12'h870:    begin Red = 8'h41;    Green = 8'h65;    Blue = 8'h8d;
end 12'h871:    begin Red = 8'h3a;    Green = 8'h60;    Blue = 8'h95;
end 12'h872:    begin Red = 8'h71;    Green = 8'h71;    Blue = 8'h4d;
end 12'h873:    begin Red = 8'h2a;    Green = 8'h55;    Blue = 8'h81;
end 12'h874:    begin Red = 8'hc7;    Green = 8'h6f;    Blue = 8'h9f;
end 12'h875:    begin Red = 8'hd5;    Green = 8'hea;    Blue = 8'hd6;
end 12'h876:    begin Red = 8'hcb;    Green = 8'h7e;    Blue = 8'ha8;
end 12'h877:    begin Red = 8'h8d;    Green = 8'hb2;    Blue = 8'h90;
end 12'h878:    begin Red = 8'h06;    Green = 8'h55;    Blue = 8'ha0;
end 12'h879:    begin Red = 8'h06;    Green = 8'h15;    Blue = 8'hff;
end 12'h87a:    begin Red = 8'h03;    Green = 8'h82;    Blue = 8'hdb;
end 12'h87b:    begin Red = 8'h5e;    Green = 8'h45;    Blue = 8'h1f;
end 12'h87c:    begin Red = 8'h6d;    Green = 8'h73;    Blue = 8'h48;
end 12'h87d:    begin Red = 8'h95;    Green = 8'hac;    Blue = 8'h81;
end 12'h87e:    begin Red = 8'h70;    Green = 8'hb0;    Blue = 8'h67;
end 12'h87f:    begin Red = 8'h71;    Green = 8'ha8;    Blue = 8'h63;
end 12'h880:    begin Red = 8'h7a;    Green = 8'h7f;    Blue = 8'h5b;
end 12'h881:    begin Red = 8'h53;    Green = 8'h85;    Blue = 8'h4a;
end 12'h882:    begin Red = 8'hf5;    Green = 8'hd3;    Blue = 8'h9d;
end 12'h883:    begin Red = 8'h83;    Green = 8'h6d;    Blue = 8'h5a;
end 12'h884:    begin Red = 8'hc4;    Green = 8'hce;    Blue = 8'ha4;
end 12'h885:    begin Red = 8'h75;    Green = 8'h6c;    Blue = 8'h5f;
end 12'h886:    begin Red = 8'ha9;    Green = 8'h50;    Blue = 8'h88;
end 12'h887:    begin Red = 8'h87;    Green = 8'h75;    Blue = 8'h59;
end 12'h888:    begin Red = 8'h04;    Green = 8'hf5;    Blue = 8'hce;
end 12'h889:    begin Red = 8'h03;    Green = 8'h82;    Blue = 8'hef;
end 12'h88a:    begin Red = 8'h02;    Green = 8'hc1;    Blue = 8'hd8;
end 12'h88b:    begin Red = 8'h58;    Green = 8'h45;    Blue = 8'h21;
end 12'h88c:    begin Red = 8'h51;    Green = 8'h3c;    Blue = 8'h23;
end 12'h88d:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'h79;
end 12'h88e:    begin Red = 8'h02;    Green = 8'h31;    Blue = 8'hd5;
end 12'h88f:    begin Red = 8'h4c;    Green = 8'h58;    Blue = 8'h3b;
end 12'h890:    begin Red = 8'ha4;    Green = 8'h51;    Blue = 8'h8d;
end 12'h891:    begin Red = 8'hd6;    Green = 8'hcc;    Blue = 8'hb3;
end 12'h892:    begin Red = 8'he0;    Green = 8'hda;    Blue = 8'hbc;
end 12'h893:    begin Red = 8'h8c;    Green = 8'ha4;    Blue = 8'h75;
end 12'h894:    begin Red = 8'h5e;    Green = 8'h4b;    Blue = 8'h25;
end 12'h895:    begin Red = 8'h52;    Green = 8'h43;    Blue = 8'h1e;
end 12'h896:    begin Red = 8'h4e;    Green = 8'h38;    Blue = 8'h19;
end 12'h897:    begin Red = 8'h02;    Green = 8'hb2;    Blue = 8'h69;
end 12'h898:    begin Red = 8'h02;    Green = 8'hd2;    Blue = 8'h8b;
end 12'h899:    begin Red = 8'h03;    Green = 8'h82;    Blue = 8'hc4;
end 12'h89a:    begin Red = 8'h90;    Green = 8'h9e;    Blue = 8'h6d;
end 12'h89b:    begin Red = 8'hbb;    Green = 8'h7a;    Blue = 8'ha9;
end 12'h89c:    begin Red = 8'h87;    Green = 8'h9c;    Blue = 8'h89;
end 12'h89d:    begin Red = 8'h47;    Green = 8'h5b;    Blue = 8'h18;
end 12'h89e:    begin Red = 8'h03;    Green = 8'hb2;    Blue = 8'hdf;
end 12'h89f:    begin Red = 8'h03;    Green = 8'hc2;    Blue = 8'hec;
end 12'h8a0:    begin Red = 8'h02;    Green = 8'h82;    Blue = 8'h1e;
end 12'h8a1:    begin Red = 8'h02;    Green = 8'ha2;    Blue = 8'h05;
end 12'h8a2:    begin Red = 8'h03;    Green = 8'h02;    Blue = 8'h9d;
end 12'h8a3:    begin Red = 8'h93;    Green = 8'hb9;    Blue = 8'h93;
end 12'h8a4:    begin Red = 8'h4d;    Green = 8'h72;    Blue = 8'h57;
end 12'h8a5:    begin Red = 8'hb4;    Green = 8'ha5;    Blue = 8'hb2;
end 12'h8a6:    begin Red = 8'h9b;    Green = 8'h4f;    Blue = 8'h86;
end 12'h8a7:    begin Red = 8'h78;    Green = 8'h66;    Blue = 8'h52;
end 12'h8a8:    begin Red = 8'h49;    Green = 8'h2e;    Blue = 8'h1f;
end 12'h8a9:    begin Red = 8'h4e;    Green = 8'h68;    Blue = 8'h17;
end 12'h8aa:    begin Red = 8'h57;    Green = 8'h34;    Blue = 8'h11;
end 12'h8ab:    begin Red = 8'h50;    Green = 8'h39;    Blue = 8'h12;
end 12'h8ac:    begin Red = 8'h76;    Green = 8'h4d;    Blue = 8'h29;
end 12'h8ad:    begin Red = 8'h63;    Green = 8'h43;    Blue = 8'h24;
end 12'h8ae:    begin Red = 8'h70;    Green = 8'h4d;    Blue = 8'h28;
end 12'h8af:    begin Red = 8'h01;    Green = 8'h91;    Blue = 8'hc9;
end 12'h8b0:    begin Red = 8'h02;    Green = 8'h72;    Blue = 8'h30;
end 12'h8b1:    begin Red = 8'ha4;    Green = 8'hae;    Blue = 8'h7c;
end 12'h8b2:    begin Red = 8'h00;    Green = 8'h18;    Blue = 8'hee;
end 12'h8b3:    begin Red = 8'h6e;    Green = 8'h66;    Blue = 8'h48;
end 12'h8b4:    begin Red = 8'hb4;    Green = 8'hb9;    Blue = 8'h8a;
end 12'h8b5:    begin Red = 8'h20;    Green = 8'h14;    Blue = 8'h17;
end 12'h8b6:    begin Red = 8'hbe;    Green = 8'hcd;    Blue = 8'hc2;
end 12'h8b7:    begin Red = 8'h65;    Green = 8'h9a;    Blue = 8'h6e;
end 12'h8b8:    begin Red = 8'he4;    Green = 8'h97;    Blue = 8'h5d;
end 12'h8b9:    begin Red = 8'he0;    Green = 8'h97;    Blue = 8'h62;
end 12'h8ba:    begin Red = 8'hdf;    Green = 8'h96;    Blue = 8'h57;
end 12'h8bb:    begin Red = 8'hfb;    Green = 8'ha1;    Blue = 8'h77;
end 12'h8bc:    begin Red = 8'hff;    Green = 8'ha2;    Blue = 8'h72;
end 12'h8bd:    begin Red = 8'h03;    Green = 8'h35;    Blue = 8'h35;
end 12'h8be:    begin Red = 8'h5e;    Green = 8'h41;    Blue = 8'h1a;
end 12'h8bf:    begin Red = 8'h04;    Green = 8'h73;    Blue = 8'h4e;
end 12'h8c0:    begin Red = 8'h65;    Green = 8'h41;    Blue = 8'h1b;
end 12'h8c1:    begin Red = 8'h9a;    Green = 8'hb0;    Blue = 8'h7c;
end 12'h8c2:    begin Red = 8'h50;    Green = 8'h37;    Blue = 8'h2c;
end 12'h8c3:    begin Red = 8'hc3;    Green = 8'hd3;    Blue = 8'ha5;
end 12'h8c4:    begin Red = 8'ha9;    Green = 8'h9e;    Blue = 8'hab;
end 12'h8c5:    begin Red = 8'hdf;    Green = 8'h96;    Blue = 8'h5d;
end 12'h8c6:    begin Red = 8'hf0;    Green = 8'h95;    Blue = 8'h67;
end 12'h8c7:    begin Red = 8'hff;    Green = 8'h9e;    Blue = 8'h6d;
end 12'h8c8:    begin Red = 8'hf8;    Green = 8'ha7;    Blue = 8'h6c;
end 12'h8c9:    begin Red = 8'h57;    Green = 8'h55;    Blue = 8'h14;
end 12'h8ca:    begin Red = 8'h74;    Green = 8'h48;    Blue = 8'h1e;
end 12'h8cb:    begin Red = 8'h4b;    Green = 8'h3b;    Blue = 8'h14;
end 12'h8cc:    begin Red = 8'h04;    Green = 8'h53;    Blue = 8'h6f;
end 12'h8cd:    begin Red = 8'h65;    Green = 8'h72;    Blue = 8'h4d;
end 12'h8ce:    begin Red = 8'h56;    Green = 8'h3a;    Blue = 8'h29;
end 12'h8cf:    begin Red = 8'h59;    Green = 8'h3a;    Blue = 8'h2f;
end 12'h8d0:    begin Red = 8'hd2;    Green = 8'hd8;    Blue = 8'ha5;
end 12'h8d1:    begin Red = 8'ha4;    Green = 8'h62;    Blue = 8'h94;
end 12'h8d2:    begin Red = 8'hbf;    Green = 8'h6d;    Blue = 8'ha0;
end 12'h8d3:    begin Red = 8'hcb;    Green = 8'hd2;    Blue = 8'hb3;
end 12'h8d4:    begin Red = 8'hff;    Green = 8'h92;    Blue = 8'h5d;
end 12'h8d5:    begin Red = 8'he6;    Green = 8'h9b;    Blue = 8'h64;
end 12'h8d6:    begin Red = 8'hcb;    Green = 8'h87;    Blue = 8'h51;
end 12'h8d7:    begin Red = 8'hc4;    Green = 8'h7f;    Blue = 8'h4c;
end 12'h8d8:    begin Red = 8'he6;    Green = 8'h91;    Blue = 8'h5a;
end 12'h8d9:    begin Red = 8'h55;    Green = 8'h3e;    Blue = 8'h19;
end 12'h8da:    begin Red = 8'h1f;    Green = 8'h30;    Blue = 8'h22;
end 12'h8db:    begin Red = 8'hac;    Green = 8'h69;    Blue = 8'h38;
end 12'h8dc:    begin Red = 8'h04;    Green = 8'hd3;    Blue = 8'h6f;
end 12'h8dd:    begin Red = 8'he1;    Green = 8'hf0;    Blue = 8'hbc;
end 12'h8de:    begin Red = 8'hc1;    Green = 8'hd0;    Blue = 8'h97;
end 12'h8df:    begin Red = 8'ha3;    Green = 8'h48;    Blue = 8'h79;
end 12'h8e0:    begin Red = 8'hd1;    Green = 8'he2;    Blue = 8'hd2;
end 12'h8e1:    begin Red = 8'hc8;    Green = 8'h76;    Blue = 8'h36;
end 12'h8e2:    begin Red = 8'hc6;    Green = 8'h71;    Blue = 8'h34;
end 12'h8e3:    begin Red = 8'hfc;    Green = 8'h9d;    Blue = 8'h63;
end 12'h8e4:    begin Red = 8'hff;    Green = 8'ha4;    Blue = 8'h66;
end 12'h8e5:    begin Red = 8'he8;    Green = 8'h8c;    Blue = 8'h4d;
end 12'h8e6:    begin Red = 8'hf7;    Green = 8'h9c;    Blue = 8'h59;
end 12'h8e7:    begin Red = 8'hf7;    Green = 8'h9c;    Blue = 8'h5f;
end 12'h8e8:    begin Red = 8'hfa;    Green = 8'ha2;    Blue = 8'h64;
end 12'h8e9:    begin Red = 8'hf0;    Green = 8'h9a;    Blue = 8'h59;
end 12'h8ea:    begin Red = 8'hf7;    Green = 8'h95;    Blue = 8'h5a;
end 12'h8eb:    begin Red = 8'hf2;    Green = 8'h93;    Blue = 8'h57;
end 12'h8ec:    begin Red = 8'he2;    Green = 8'h88;    Blue = 8'h48;
end 12'h8ed:    begin Red = 8'hd5;    Green = 8'h80;    Blue = 8'h43;
end 12'h8ee:    begin Red = 8'hfe;    Green = 8'h94;    Blue = 8'h4a;
end 12'h8ef:    begin Red = 8'hc2;    Green = 8'h7a;    Blue = 8'h45;
end 12'h8f0:    begin Red = 8'hec;    Green = 8'h95;    Blue = 8'h5d;
end 12'h8f1:    begin Red = 8'hf5;    Green = 8'ha1;    Blue = 8'h67;
end 12'h8f2:    begin Red = 8'h50;    Green = 8'h40;    Blue = 8'h19;
end 12'h8f3:    begin Red = 8'h21;    Green = 8'h2e;    Blue = 8'h1d;
end 12'h8f4:    begin Red = 8'hb9;    Green = 8'h71;    Blue = 8'h3c;
end 12'h8f5:    begin Red = 8'hcb;    Green = 8'h72;    Blue = 8'h43;
end 12'h8f6:    begin Red = 8'hd5;    Green = 8'h7a;    Blue = 8'h45;
end 12'h8f7:    begin Red = 8'had;    Green = 8'hc5;    Blue = 8'h92;
end 12'h8f8:    begin Red = 8'had;    Green = 8'ha9;    Blue = 8'h7e;
end 12'h8f9:    begin Red = 8'ha4;    Green = 8'h90;    Blue = 8'h6a;
end 12'h8fa:    begin Red = 8'h9e;    Green = 8'h61;    Blue = 8'h91;
end 12'h8fb:    begin Red = 8'h9e;    Green = 8'h49;    Blue = 8'h83;
end 12'h8fc:    begin Red = 8'he3;    Green = 8'h9d;    Blue = 8'h55;
end 12'h8fd:    begin Red = 8'h73;    Green = 8'h9f;    Blue = 8'h80;
end 12'h8fe:    begin Red = 8'h1f;    Green = 8'h2d;    Blue = 8'h18;
end 12'h8ff:    begin Red = 8'h53;    Green = 8'h45;    Blue = 8'h25;
end 12'h900:    begin Red = 8'h02;    Green = 8'hf2;    Blue = 8'h99;
end 12'h901:    begin Red = 8'hb0;    Green = 8'hc4;    Blue = 8'h9d;
end 12'h902:    begin Red = 8'h7d;    Green = 8'h77;    Blue = 8'h4f;
end 12'h903:    begin Red = 8'hfc;    Green = 8'hdd;    Blue = 8'ha1;
end 12'h904:    begin Red = 8'hf4;    Green = 8'hde;    Blue = 8'h9c;
end 12'h905:    begin Red = 8'hff;    Green = 8'hdf;    Blue = 8'h9c;
end 12'h906:    begin Red = 8'h49;    Green = 8'h2f;    Blue = 8'h28;
end 12'h907:    begin Red = 8'hdf;    Green = 8'hb7;    Blue = 8'h90;
end 12'h908:    begin Red = 8'h99;    Green = 8'h44;    Blue = 8'h7f;
end 12'h909:    begin Red = 8'hdc;    Green = 8'h97;    Blue = 8'h68;
end 12'h90a:    begin Red = 8'hea;    Green = 8'h93;    Blue = 8'h6c;
end 12'h90b:    begin Red = 8'h65;    Green = 8'ha6;    Blue = 8'h81;
end 12'h90c:    begin Red = 8'hc4;    Green = 8'h8d;    Blue = 8'h56;
end 12'h90d:    begin Red = 8'hcc;    Green = 8'h8e;    Blue = 8'h57;
end 12'h90e:    begin Red = 8'hca;    Green = 8'h79;    Blue = 8'h3b;
end 12'h90f:    begin Red = 8'hb3;    Green = 8'h6f;    Blue = 8'h3a;
end 12'h910:    begin Red = 8'hb5;    Green = 8'h6a;    Blue = 8'h38;
end 12'h911:    begin Red = 8'hce;    Green = 8'he0;    Blue = 8'hb9;
end 12'h912:    begin Red = 8'h8f;    Green = 8'h97;    Blue = 8'h72;
end 12'h913:    begin Red = 8'h82;    Green = 8'h96;    Blue = 8'h7f;
end 12'h914:    begin Red = 8'hbd;    Green = 8'h69;    Blue = 8'h3c;
end 12'h915:    begin Red = 8'h35;    Green = 8'h26;    Blue = 8'h22;
end 12'h916:    begin Red = 8'hf4;    Green = 8'hd8;    Blue = 8'ha3;
end 12'h917:    begin Red = 8'hd9;    Green = 8'h9f;    Blue = 8'h61;
end 12'h918:    begin Red = 8'hdf;    Green = 8'h9c;    Blue = 8'h64;
end 12'h919:    begin Red = 8'h5b;    Green = 8'ha6;    Blue = 8'h81;
end 12'h91a:    begin Red = 8'h71;    Green = 8'ha0;    Blue = 8'h87;
end 12'h91b:    begin Red = 8'hee;    Green = 8'h90;    Blue = 8'h67;
end 12'h91c:    begin Red = 8'hcb;    Green = 8'h94;    Blue = 8'h5d;
end 12'h91d:    begin Red = 8'hd9;    Green = 8'h94;    Blue = 8'h5f;
end 12'h91e:    begin Red = 8'h35;    Green = 8'h40;    Blue = 8'h2a;
end 12'h91f:    begin Red = 8'h0d;    Green = 8'h26;    Blue = 8'h12;
end 12'h920:    begin Red = 8'hbe;    Green = 8'h6f;    Blue = 8'h30;
end 12'h921:    begin Red = 8'hd3;    Green = 8'he4;    Blue = 8'hbd;
end 12'h922:    begin Red = 8'h78;    Green = 8'hab;    Blue = 8'h8a;
end 12'h923:    begin Red = 8'h89;    Green = 8'h98;    Blue = 8'h69;
end 12'h924:    begin Red = 8'h8c;    Green = 8'h45;    Blue = 8'h78;
end 12'h925:    begin Red = 8'h8d;    Green = 8'h9c;    Blue = 8'h7a;
end 12'h926:    begin Red = 8'ha9;    Green = 8'h6e;    Blue = 8'h3b;
end 12'h927:    begin Red = 8'hab;    Green = 8'hbf;    Blue = 8'h96;
end 12'h928:    begin Red = 8'hc6;    Green = 8'h60;    Blue = 8'h1a;
end 12'h929:    begin Red = 8'h74;    Green = 8'hbe;    Blue = 8'hd1;
end 12'h92a:    begin Red = 8'h69;    Green = 8'hce;    Blue = 8'he9;
end 12'h92b:    begin Red = 8'h35;    Green = 8'h53;    Blue = 8'h86;
end 12'h92c:    begin Red = 8'h78;    Green = 8'h91;    Blue = 8'hf4;
end 12'h92d:    begin Red = 8'h35;    Green = 8'h4e;    Blue = 8'h94;
end 12'h92e:    begin Red = 8'h7b;    Green = 8'h9b;    Blue = 8'hf6;
end 12'h92f:    begin Red = 8'h7a;    Green = 8'h5d;    Blue = 8'h4f;
end 12'h930:    begin Red = 8'h9b;    Green = 8'h5c;    Blue = 8'h8b;
end 12'h931:    begin Red = 8'h90;    Green = 8'h55;    Blue = 8'h84;
end 12'h932:    begin Red = 8'ha9;    Green = 8'h5f;    Blue = 8'h93;
end 12'h933:    begin Red = 8'ha2;    Green = 8'h59;    Blue = 8'h94;
end 12'h934:    begin Red = 8'had;    Green = 8'h46;    Blue = 8'h8c;
end 12'h935:    begin Red = 8'h6a;    Green = 8'hae;    Blue = 8'h89;
end 12'h936:    begin Red = 8'hde;    Green = 8'h91;    Blue = 8'h59;
end 12'h937:    begin Red = 8'hb0;    Green = 8'h61;    Blue = 8'h2f;
end 12'h938:    begin Red = 8'hbd;    Green = 8'h67;    Blue = 8'h2f;
end 12'h939:    begin Red = 8'hc8;    Green = 8'h5f;    Blue = 8'h20;
end 12'h93a:    begin Red = 8'h6c;    Green = 8'hca;    Blue = 8'hee;
end 12'h93b:    begin Red = 8'h36;    Green = 8'h55;    Blue = 8'h8c;
end 12'h93c:    begin Red = 8'h40;    Green = 8'h4e;    Blue = 8'h85;
end 12'h93d:    begin Red = 8'h3e;    Green = 8'h51;    Blue = 8'h8c;
end 12'h93e:    begin Red = 8'h6e;    Green = 8'ha3;    Blue = 8'hf6;
end 12'h93f:    begin Red = 8'h37;    Green = 8'h58;    Blue = 8'h91;
end 12'h940:    begin Red = 8'h66;    Green = 8'h9c;    Blue = 8'he9;
end 12'h941:    begin Red = 8'haa;    Green = 8'hac;    Blue = 8'hb3;
end 12'h942:    begin Red = 8'h96;    Green = 8'h48;    Blue = 8'h88;
end 12'h943:    begin Red = 8'h91;    Green = 8'h40;    Blue = 8'h7a;
end 12'h944:    begin Red = 8'hab;    Green = 8'h5a;    Blue = 8'h93;
end 12'h945:    begin Red = 8'h9e;    Green = 8'h4e;    Blue = 8'h8c;
end 12'h946:    begin Red = 8'hef;    Green = 8'ha1;    Blue = 8'h6b;
end 12'h947:    begin Red = 8'h5b;    Green = 8'ha7;    Blue = 8'h8c;
end 12'h948:    begin Red = 8'h6a;    Green = 8'ha1;    Blue = 8'h7f;
end 12'h949:    begin Red = 8'he2;    Green = 8'h9c;    Blue = 8'h5e;
end 12'h94a:    begin Red = 8'hbf;    Green = 8'h77;    Blue = 8'h40;
end 12'h94b:    begin Red = 8'hae;    Green = 8'h67;    Blue = 8'h32;
end 12'h94c:    begin Red = 8'h8c;    Green = 8'h8f;    Blue = 8'h65;
end 12'h94d:    begin Red = 8'hb6;    Green = 8'h65;    Blue = 8'h31;
end 12'h94e:    begin Red = 8'h50;    Green = 8'hdf;    Blue = 8'hf6;
end 12'h94f:    begin Red = 8'h5b;    Green = 8'hcd;    Blue = 8'hee;
end 12'h950:    begin Red = 8'h59;    Green = 8'hc8;    Blue = 8'hea;
end 12'h951:    begin Red = 8'h61;    Green = 8'hca;    Blue = 8'hee;
end 12'h952:    begin Red = 8'h60;    Green = 8'hd7;    Blue = 8'hf6;
end 12'h953:    begin Red = 8'he6;    Green = 8'h90;    Blue = 8'h63;
end 12'h954:    begin Red = 8'h76;    Green = 8'h9e;    Blue = 8'h87;
end 12'h955:    begin Red = 8'hdd;    Green = 8'h95;    Blue = 8'h4f;
end 12'h956:    begin Red = 8'hc4;    Green = 8'hd8;    Blue = 8'hb0;
end 12'h957:    begin Red = 8'hd0;    Green = 8'h82;    Blue = 8'h4c;
end 12'h958:    begin Red = 8'hbf;    Green = 8'h7b;    Blue = 8'h4e;
end 12'h959:    begin Red = 8'hbc;    Green = 8'h76;    Blue = 8'h4d;
end 12'h95a:    begin Red = 8'hca;    Green = 8'h84;    Blue = 8'h4b;
end 12'h95b:    begin Red = 8'hd3;    Green = 8'h88;    Blue = 8'h52;
end 12'h95c:    begin Red = 8'hc3;    Green = 8'h98;    Blue = 8'h61;
end 12'h95d:    begin Red = 8'hb9;    Green = 8'h8e;    Blue = 8'h61;
end 12'h95e:    begin Red = 8'h7c;    Green = 8'h71;    Blue = 8'h4b;
end 12'h95f:    begin Red = 8'h9f;    Green = 8'had;    Blue = 8'ha9;
end 12'h960:    begin Red = 8'h5f;    Green = 8'ha8;    Blue = 8'h87;
end 12'h961:    begin Red = 8'he0;    Green = 8'ha5;    Blue = 8'h5f;
end 12'h962:    begin Red = 8'hc7;    Green = 8'h7d;    Blue = 8'h47;
end 12'h963:    begin Red = 8'hee;    Green = 8'h9f;    Blue = 8'h65;
end 12'h964:    begin Red = 8'hbf;    Green = 8'h72;    Blue = 8'h3d;
end 12'h965:    begin Red = 8'hb8;    Green = 8'h7b;    Blue = 8'h54;
end 12'h966:    begin Red = 8'hce;    Green = 8'h7e;    Blue = 8'h44;
end 12'h967:    begin Red = 8'hcb;    Green = 8'h93;    Blue = 8'h6d;
end 12'h968:    begin Red = 8'hcd;    Green = 8'hd8;    Blue = 8'ha9;
end 12'h969:    begin Red = 8'hc0;    Green = 8'h95;    Blue = 8'h56;
end 12'h96a:    begin Red = 8'hd4;    Green = 8'hdc;    Blue = 8'hbe;
end 12'h96b:    begin Red = 8'ha6;    Green = 8'h6c;    Blue = 8'h95;
end 12'h96c:    begin Red = 8'hcb;    Green = 8'h81;    Blue = 8'h54;
end 12'h96d:    begin Red = 8'hca;    Green = 8'h84;    Blue = 8'h59;
end 12'h96e:    begin Red = 8'hbe;    Green = 8'h80;    Blue = 8'h52;
end 12'h96f:    begin Red = 8'hc1;    Green = 8'h7e;    Blue = 8'h5a;
end 12'h970:    begin Red = 8'ha4;    Green = 8'h63;    Blue = 8'h32;
end 12'h971:    begin Red = 8'h84;    Green = 8'h95;    Blue = 8'h73;
end 12'h972:    begin Red = 8'heb;    Green = 8'h9f;    Blue = 8'h5f;
end 12'h973:    begin Red = 8'hc1;    Green = 8'h85;    Blue = 8'hae;
end 12'h974:    begin Red = 8'hac;    Green = 8'h74;    Blue = 8'h9a;
end 12'h975:    begin Red = 8'hc6;    Green = 8'h8b;    Blue = 8'hb4;
end 12'h976:    begin Red = 8'hc6;    Green = 8'h86;    Blue = 8'hb0;
end 12'h977:    begin Red = 8'h87;    Green = 8'h59;    Blue = 8'h77;
end 12'h978:    begin Red = 8'h97;    Green = 8'h66;    Blue = 8'h8c;
end 12'h979:    begin Red = 8'h9d;    Green = 8'h6d;    Blue = 8'h8d;
end 12'h97a:    begin Red = 8'h8d;    Green = 8'h90;    Blue = 8'h6e;
end 12'h97b:    begin Red = 8'hb0;    Green = 8'h9f;    Blue = 8'ha2;
end 12'h97c:    begin Red = 8'ha3;    Green = 8'h53;    Blue = 8'h7f;
end 12'h97d:    begin Red = 8'h9d;    Green = 8'h55;    Blue = 8'h8d;
end 12'h97e:    begin Red = 8'h6a;    Green = 8'h66;    Blue = 8'h6a;
end 12'h97f:    begin Red = 8'h72;    Green = 8'h6f;    Blue = 8'h6d;
end 12'h980:    begin Red = 8'h73;    Green = 8'h6e;    Blue = 8'h7a;
end 12'h981:    begin Red = 8'ha3;    Green = 8'h94;    Blue = 8'h7f;
end 12'h982:    begin Red = 8'ha8;    Green = 8'h93;    Blue = 8'h81;
end 12'h983:    begin Red = 8'h71;    Green = 8'h71;    Blue = 8'h68;
end 12'h984:    begin Red = 8'haa;    Green = 8'h96;    Blue = 8'h87;
end 12'h985:    begin Red = 8'h5a;    Green = 8'h5a;    Blue = 8'h5a;
end 12'h986:    begin Red = 8'hcb;    Green = 8'he0;    Blue = 8'hb2;
end 12'h987:    begin Red = 8'hb7;    Green = 8'h79;    Blue = 8'ha0;
end 12'h988:    begin Red = 8'hb1;    Green = 8'h75;    Blue = 8'h9d;
end 12'h989:    begin Red = 8'h9e;    Green = 8'h68;    Blue = 8'h8e;
end 12'h98a:    begin Red = 8'h9b;    Green = 8'h41;    Blue = 8'h8f;
end 12'h98b:    begin Red = 8'h93;    Green = 8'h43;    Blue = 8'h81;
end 12'h98c:    begin Red = 8'hea;    Green = 8'h96;    Blue = 8'h65;
end 12'h98d:    begin Red = 8'h5c;    Green = 8'had;    Blue = 8'h90;
end 12'h98e:    begin Red = 8'h66;    Green = 8'h6f;    Blue = 8'h6e;
end 12'h98f:    begin Red = 8'hb8;    Green = 8'ha0;    Blue = 8'h85;
end 12'h990:    begin Red = 8'h6a;    Green = 8'h6c;    Blue = 8'h7a;
end 12'h991:    begin Red = 8'h74;    Green = 8'h76;    Blue = 8'h78;
end 12'h992:    begin Red = 8'hc3;    Green = 8'ha9;    Blue = 8'h8c;
end 12'h993:    begin Red = 8'h6b;    Green = 8'h6d;    Blue = 8'h73;
end 12'h994:    begin Red = 8'hbd;    Green = 8'ha8;    Blue = 8'h85;
end 12'h995:    begin Red = 8'h70;    Green = 8'h68;    Blue = 8'h77;
end 12'h996:    begin Red = 8'h61;    Green = 8'h6a;    Blue = 8'h73;
end 12'h997:    begin Red = 8'h64;    Green = 8'h70;    Blue = 8'h76;
end 12'h998:    begin Red = 8'h5c;    Green = 8'h5e;    Blue = 8'h61;
end 12'h999:    begin Red = 8'h89;    Green = 8'h98;    Blue = 8'h74;
end 12'h99a:    begin Red = 8'h62;    Green = 8'h96;    Blue = 8'h57;
end 12'h99b:    begin Red = 8'h61;    Green = 8'h93;    Blue = 8'h52;
end 12'h99c:    begin Red = 8'h88;    Green = 8'h59;    Blue = 8'h7d;
end 12'h99d:    begin Red = 8'h9b;    Green = 8'h61;    Blue = 8'h86;
end 12'h99e:    begin Red = 8'hcd;    Green = 8'hc2;    Blue = 8'hc2;
end 12'h99f:    begin Red = 8'ha9;    Green = 8'h61;    Blue = 8'h2b;
end 12'h9a0:    begin Red = 8'h65;    Green = 8'h41;    Blue = 8'h3a;
end 12'h9a1:    begin Red = 8'h8f;    Green = 8'h82;    Blue = 8'h58;
end 12'h9a2:    begin Red = 8'h93;    Green = 8'h85;    Blue = 8'h61;
end 12'h9a3:    begin Red = 8'h8a;    Green = 8'h7c;    Blue = 8'h58;
end 12'h9a4:    begin Red = 8'h9e;    Green = 8'h63;    Blue = 8'h3c;
end 12'h9a5:    begin Red = 8'ha5;    Green = 8'hb8;    Blue = 8'h94;
end 12'h9a6:    begin Red = 8'h85;    Green = 8'h54;    Blue = 8'h77;
end 12'h9a7:    begin Red = 8'hb2;    Green = 8'haa;    Blue = 8'hb2;
end 12'h9a8:    begin Red = 8'ha9;    Green = 8'hb8;    Blue = 8'hae;
end 12'h9a9:    begin Red = 8'h9b;    Green = 8'h52;    Blue = 8'h81;
end 12'h9aa:    begin Red = 8'h75;    Green = 8'hb3;    Blue = 8'h95;
end 12'h9ab:    begin Red = 8'h72;    Green = 8'ha7;    Blue = 8'h87;
end 12'h9ac:    begin Red = 8'h7c;    Green = 8'hae;    Blue = 8'h85;
end 12'h9ad:    begin Red = 8'h89;    Green = 8'hb1;    Blue = 8'h8a;
end 12'h9ae:    begin Red = 8'h5d;    Green = 8'h4d;    Blue = 8'h48;
end 12'h9af:    begin Red = 8'h90;    Green = 8'h87;    Blue = 8'h57;
end 12'h9b0:    begin Red = 8'h7c;    Green = 8'h7f;    Blue = 8'h4b;
end 12'h9b1:    begin Red = 8'h93;    Green = 8'h61;    Blue = 8'h42;
end 12'h9b2:    begin Red = 8'hbb;    Green = 8'h75;    Blue = 8'h52;
end 12'h9b3:    begin Red = 8'ha3;    Green = 8'h61;    Blue = 8'h9d;
end 12'h9b4:    begin Red = 8'h5a;    Green = 8'h48;    Blue = 8'h3d;
end 12'h9b5:    begin Red = 8'hd3;    Green = 8'h87;    Blue = 8'h64;
end 12'h9b6:    begin Red = 8'haa;    Green = 8'hca;    Blue = 8'ha1;
end 12'h9b7:    begin Red = 8'h99;    Green = 8'h66;    Blue = 8'h42;
end 12'h9b8:    begin Red = 8'hed;    Green = 8'hcd;    Blue = 8'ha5;
end 12'h9b9:    begin Red = 8'h95;    Green = 8'h57;    Blue = 8'h7e;
end 12'h9ba:    begin Red = 8'h8d;    Green = 8'h30;    Blue = 8'h70;
end 12'h9bb:    begin Red = 8'hba;    Green = 8'h9a;    Blue = 8'h66;
end 12'h9bc:    begin Red = 8'haf;    Green = 8'h98;    Blue = 8'h67;
end 12'h9bd:    begin Red = 8'h95;    Green = 8'h92;    Blue = 8'h63;
end 12'h9be:    begin Red = 8'h4d;    Green = 8'h45;    Blue = 8'h3e;
end 12'h9bf:    begin Red = 8'hde;    Green = 8'he9;    Blue = 8'hb1;
end 12'h9c0:    begin Red = 8'ha2;    Green = 8'haa;    Blue = 8'h82;
end 12'h9c1:    begin Red = 8'had;    Green = 8'hb1;    Blue = 8'hbc;
end 12'h9c2:    begin Red = 8'hb9;    Green = 8'hc3;    Blue = 8'hb1;
end 12'h9c3:    begin Red = 8'hb0;    Green = 8'hc1;    Blue = 8'ha7;
end 12'h9c4:    begin Red = 8'h98;    Green = 8'h4c;    Blue = 8'h81;
end 12'h9c5:    begin Red = 8'h98;    Green = 8'h35;    Blue = 8'h6d;
end 12'h9c6:    begin Red = 8'h84;    Green = 8'hb0;    Blue = 8'h89;
end 12'h9c7:    begin Red = 8'h72;    Green = 8'haa;    Blue = 8'h75;
end 12'h9c8:    begin Red = 8'hc8;    Green = 8'hc0;    Blue = 8'ha4;
end 12'h9c9:    begin Red = 8'hcb;    Green = 8'hc4;    Blue = 8'haa;
end 12'h9ca:    begin Red = 8'hd7;    Green = 8'hdc;    Blue = 8'ha4;
end 12'h9cb:    begin Red = 8'hc8;    Green = 8'hc6;    Blue = 8'h9d;
end 12'h9cc:    begin Red = 8'h9a;    Green = 8'h60;    Blue = 8'h42;
end 12'h9cd:    begin Red = 8'ha8;    Green = 8'h9f;    Blue = 8'h71;
end 12'h9ce:    begin Red = 8'ha6;    Green = 8'h8f;    Blue = 8'h63;
end 12'h9cf:    begin Red = 8'ha9;    Green = 8'h69;    Blue = 8'h9a;
end 12'h9d0:    begin Red = 8'ha4;    Green = 8'h62;    Blue = 8'h81;
end 12'h9d1:    begin Red = 8'hef;    Green = 8'hd7;    Blue = 8'hba;
end 12'h9d2:    begin Red = 8'hc3;    Green = 8'hb5;    Blue = 8'h98;
end 12'h9d3:    begin Red = 8'h98;    Green = 8'h99;    Blue = 8'h78;
end 12'h9d4:    begin Red = 8'h92;    Green = 8'h99;    Blue = 8'h7a;
end 12'h9d5:    begin Red = 8'h90;    Green = 8'h70;    Blue = 8'h36;
end 12'h9d6:    begin Red = 8'h45;    Green = 8'h54;    Blue = 8'h81;
end 12'h9d7:    begin Red = 8'h75;    Green = 8'ha1;    Blue = 8'he8;
end 12'h9d8:    begin Red = 8'h7a;    Green = 8'h4c;    Blue = 8'h74;
end 12'h9d9:    begin Red = 8'h7b;    Green = 8'h4c;    Blue = 8'h6d;
end 12'h9da:    begin Red = 8'h6c;    Green = 8'h3d;    Blue = 8'h5f;
end 12'h9db:    begin Red = 8'h68;    Green = 8'h49;    Blue = 8'h61;
end 12'h9dc:    begin Red = 8'h74;    Green = 8'h4b;    Blue = 8'h6d;
end 12'h9dd:    begin Red = 8'h6f;    Green = 8'h42;    Blue = 8'h63;
end 12'h9de:    begin Red = 8'h77;    Green = 8'h46;    Blue = 8'h69;
end 12'h9df:    begin Red = 8'hc3;    Green = 8'hcd;    Blue = 8'h9c;
end 12'h9e0:    begin Red = 8'h3a;    Green = 8'h5b;    Blue = 8'h7e;
end 12'h9e1:    begin Red = 8'h74;    Green = 8'h94;    Blue = 8'hef;
end 12'h9e2:    begin Red = 8'h81;    Green = 8'h65;    Blue = 8'h37;
end 12'h9e3:    begin Red = 8'hff;    Green = 8'hed;    Blue = 8'hcc;
end 12'h9e4:    begin Red = 8'hef;    Green = 8'hdf;    Blue = 8'hbd;
end 12'h9e5:    begin Red = 8'hdc;    Green = 8'hcf;    Blue = 8'haf;
end 12'h9e6:    begin Red = 8'h6d;    Green = 8'h5c;    Blue = 8'h44;
end 12'h9e7:    begin Red = 8'hbb;    Green = 8'hab;    Blue = 8'h8d;
end 12'h9e8:    begin Red = 8'hdc;    Green = 8'hd5;    Blue = 8'hb4;
end 12'h9e9:    begin Red = 8'haf;    Green = 8'ha4;    Blue = 8'h90;
end 12'h9ea:    begin Red = 8'hb8;    Green = 8'hae;    Blue = 8'h96;
end 12'h9eb:    begin Red = 8'hee;    Green = 8'he7;    Blue = 8'hc8;
end 12'h9ec:    begin Red = 8'h79;    Green = 8'ha6;    Blue = 8'hf6;
end 12'h9ed:    begin Red = 8'h6f;    Green = 8'h98;    Blue = 8'hf1;
end 12'h9ee:    begin Red = 8'h74;    Green = 8'h9d;    Blue = 8'hf6;
end 12'h9ef:    begin Red = 8'h66;    Green = 8'h33;    Blue = 8'h6f;
end 12'h9f0:    begin Red = 8'h62;    Green = 8'h2e;    Blue = 8'h64;
end 12'h9f1:    begin Red = 8'h57;    Green = 8'h26;    Blue = 8'h5b;
end 12'h9f2:    begin Red = 8'h5a;    Green = 8'h21;    Blue = 8'h55;
end 12'h9f3:    begin Red = 8'h6d;    Green = 8'h35;    Blue = 8'h73;
end 12'h9f4:    begin Red = 8'h6e;    Green = 8'h38;    Blue = 8'h6b;
end 12'h9f5:    begin Red = 8'h6b;    Green = 8'h33;    Blue = 8'h67;
end 12'h9f6:    begin Red = 8'h5f;    Green = 8'h2d;    Blue = 8'h5f;
end 12'h9f7:    begin Red = 8'h72;    Green = 8'h34;    Blue = 8'h74;
end 12'h9f8:    begin Red = 8'h77;    Green = 8'h96;    Blue = 8'hf6;
end 12'h9f9:    begin Red = 8'hd6;    Green = 8'heb;    Blue = 8'hd1;
end 12'h9fa:    begin Red = 8'h60;    Green = 8'h59;    Blue = 8'h42;
end 12'h9fb:    begin Red = 8'hc8;    Green = 8'hba;    Blue = 8'h9d;
end 12'h9fc:    begin Red = 8'h98;    Green = 8'h81;    Blue = 8'h66;
end 12'h9fd:    begin Red = 8'he6;    Green = 8'hd9;    Blue = 8'hb9;
end 12'h9fe:    begin Red = 8'hca;    Green = 8'hd1;    Blue = 8'h9e;
end 12'h9ff:    begin Red = 8'he4;    Green = 8'he1;    Blue = 8'h9b;
end 12'ha00:    begin Red = 8'hd7;    Green = 8'hb7;    Blue = 8'h7f;
end 12'ha01:    begin Red = 8'haf;    Green = 8'h98;    Blue = 8'h79;
end 12'ha02:    begin Red = 8'h5b;    Green = 8'h50;    Blue = 8'h4d;
end 12'ha03:    begin Red = 8'h8d;    Green = 8'h52;    Blue = 8'h75;
end 12'ha04:    begin Red = 8'h9a;    Green = 8'h49;    Blue = 8'h7b;
end 12'ha05:    begin Red = 8'hcd;    Green = 8'hbd;    Blue = 8'h9f;
end 12'ha06:    begin Red = 8'ha1;    Green = 8'ha0;    Blue = 8'h7e;
end 12'ha07:    begin Red = 8'h01;    Green = 8'h8f;    Blue = 8'h13;
end 12'ha08:    begin Red = 8'h64;    Green = 8'h4e;    Blue = 8'h3c;
end 12'ha09:    begin Red = 8'h38;    Green = 8'h53;    Blue = 8'h75;
end 12'ha0a:    begin Red = 8'ha9;    Green = 8'h97;    Blue = 8'h63;
end 12'ha0b:    begin Red = 8'ha2;    Green = 8'h7f;    Blue = 8'h58;
end 12'ha0c:    begin Red = 8'h93;    Green = 8'h8f;    Blue = 8'h97;
end 12'ha0d:    begin Red = 8'h9c;    Green = 8'h8c;    Blue = 8'h98;
end 12'ha0e:    begin Red = 8'hea;    Green = 8'hde;    Blue = 8'hc0;
end 12'ha0f:    begin Red = 8'hec;    Green = 8'hdd;    Blue = 8'hc5;
end 12'ha10:    begin Red = 8'hdc;    Green = 8'hd1;    Blue = 8'hbb;
end 12'ha11:    begin Red = 8'hf2;    Green = 8'hee;    Blue = 8'hd5;
end 12'ha12:    begin Red = 8'hbd;    Green = 8'hb7;    Blue = 8'h9b;
end 12'ha13:    begin Red = 8'h52;    Green = 8'h36;    Blue = 8'h23;
end 12'ha14:    begin Red = 8'he4;    Green = 8'hb6;    Blue = 8'h86;
end 12'ha15:    begin Red = 8'h2d;    Green = 8'h56;    Blue = 8'h8e;
end 12'ha16:    begin Red = 8'hb4;    Green = 8'h96;    Blue = 8'h63;
end 12'ha17:    begin Red = 8'h97;    Green = 8'h79;    Blue = 8'h4b;
end 12'ha18:    begin Red = 8'hcc;    Green = 8'hcb;    Blue = 8'ha7;
end 12'ha19:    begin Red = 8'he6;    Green = 8'hd4;    Blue = 8'h93;
end 12'ha1a:    begin Red = 8'h8e;    Green = 8'h68;    Blue = 8'h53;
end 12'ha1b:    begin Red = 8'ha7;    Green = 8'ha4;    Blue = 8'ha5;
end 12'ha1c:    begin Red = 8'hff;    Green = 8'hf5;    Blue = 8'he6;
end 12'ha1d:    begin Red = 8'hfc;    Green = 8'hf3;    Blue = 8'he0;
end 12'ha1e:    begin Red = 8'hfb;    Green = 8'hf0;    Blue = 8'hd7;
end 12'ha1f:    begin Red = 8'hfc;    Green = 8'hfc;    Blue = 8'he2;
end 12'ha20:    begin Red = 8'hfb;    Green = 8'hf7;    Blue = 8'hd7;
end 12'ha21:    begin Red = 8'hf5;    Green = 8'he6;    Blue = 8'hca;
end 12'ha22:    begin Red = 8'h7b;    Green = 8'h7e;    Blue = 8'h83;
end 12'ha23:    begin Red = 8'h7a;    Green = 8'h7d;    Blue = 8'h7d;
end 12'ha24:    begin Red = 8'haf;    Green = 8'hb9;    Blue = 8'h86;
end 12'ha25:    begin Red = 8'h5e;    Green = 8'h3c;    Blue = 8'h2c;
end 12'ha26:    begin Red = 8'h73;    Green = 8'h68;    Blue = 8'h5a;
end 12'ha27:    begin Red = 8'h9e;    Green = 8'h92;    Blue = 8'h85;
end 12'ha28:    begin Red = 8'ha5;    Green = 8'h90;    Blue = 8'h86;
end 12'ha29:    begin Red = 8'h85;    Green = 8'h6e;    Blue = 8'h3b;
end 12'ha2a:    begin Red = 8'he4;    Green = 8'he0;    Blue = 8'hb3;
end 12'ha2b:    begin Red = 8'h86;    Green = 8'h6c;    Blue = 8'h35;
end 12'ha2c:    begin Red = 8'hd4;    Green = 8'hc3;    Blue = 8'h7e;
end 12'ha2d:    begin Red = 8'hd7;    Green = 8'hbc;    Blue = 8'h7a;
end 12'ha2e:    begin Red = 8'hf7;    Green = 8'hee;    Blue = 8'hd2;
end 12'ha2f:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h3f;
end 12'ha30:    begin Red = 8'he1;    Green = 8'hbe;    Blue = 8'h8e;
end 12'ha31:    begin Red = 8'hb4;    Green = 8'ha8;    Blue = 8'h9b;
end 12'ha32:    begin Red = 8'haf;    Green = 8'h79;    Blue = 8'h55;
end 12'ha33:    begin Red = 8'haf;    Green = 8'h72;    Blue = 8'h35;
end 12'ha34:    begin Red = 8'he3;    Green = 8'hc0;    Blue = 8'h94;
end 12'ha35:    begin Red = 8'ha0;    Green = 8'h9a;    Blue = 8'h98;
end 12'ha36:    begin Red = 8'h07;    Green = 8'h05;    Blue = 8'hac;
end 12'ha37:    begin Red = 8'hf2;    Green = 8'hdf;    Blue = 8'hc6;
end 12'ha38:    begin Red = 8'he5;    Green = 8'hda;    Blue = 8'hc3;
end 12'ha39:    begin Red = 8'h73;    Green = 8'h5c;    Blue = 8'h13;
end 12'ha3a:    begin Red = 8'heb;    Green = 8'he1;    Blue = 8'hcd;
end 12'ha3b:    begin Red = 8'he2;    Green = 8'hd3;    Blue = 8'hbe;
end 12'ha3c:    begin Red = 8'hb0;    Green = 8'ha9;    Blue = 8'h93;
end 12'ha3d:    begin Red = 8'hb7;    Green = 8'ha5;    Blue = 8'hab;
end 12'ha3e:    begin Red = 8'h7e;    Green = 8'h6e;    Blue = 8'h36;
end 12'ha3f:    begin Red = 8'h70;    Green = 8'h50;    Blue = 8'h17;
end 12'ha40:    begin Red = 8'h7f;    Green = 8'h6c;    Blue = 8'h3d;
end 12'ha41:    begin Red = 8'h69;    Green = 8'h55;    Blue = 8'h10;
end 12'ha42:    begin Red = 8'hf2;    Green = 8'he0;    Blue = 8'hcb;
end 12'ha43:    begin Red = 8'ha8;    Green = 8'h9a;    Blue = 8'h7e;
end 12'ha44:    begin Red = 8'h60;    Green = 8'h90;    Blue = 8'h68;
end 12'ha45:    begin Red = 8'hae;    Green = 8'hb9;    Blue = 8'h81;
end 12'ha46:    begin Red = 8'hb3;    Green = 8'ha2;    Blue = 8'h88;
end 12'ha47:    begin Red = 8'hbd;    Green = 8'hbf;    Blue = 8'haa;
end 12'ha48:    begin Red = 8'hcc;    Green = 8'hb4;    Blue = 8'ha3;
end 12'ha49:    begin Red = 8'hca;    Green = 8'hbb;    Blue = 8'ha7;
end 12'ha4a:    begin Red = 8'hc8;    Green = 8'hb7;    Blue = 8'hb0;
end 12'ha4b:    begin Red = 8'hd5;    Green = 8'hc3;    Blue = 8'hb2;
end 12'ha4c:    begin Red = 8'hc4;    Green = 8'hb6;    Blue = 8'ha4;
end 12'ha4d:    begin Red = 8'h87;    Green = 8'h6e;    Blue = 8'h2f;
end 12'ha4e:    begin Red = 8'hee;    Green = 8'hda;    Blue = 8'hcb;
end 12'ha4f:    begin Red = 8'h72;    Green = 8'h5c;    Blue = 8'h1b;
end 12'ha50:    begin Red = 8'hfb;    Green = 8'hf8;    Blue = 8'heb;
end 12'ha51:    begin Red = 8'hb3;    Green = 8'ha3;    Blue = 8'h95;
end 12'ha52:    begin Red = 8'ha8;    Green = 8'hb3;    Blue = 8'h94;
end 12'ha53:    begin Red = 8'h9b;    Green = 8'h6e;    Blue = 8'h27;
end 12'ha54:    begin Red = 8'h95;    Green = 8'h9d;    Blue = 8'ha2;
end 12'ha55:    begin Red = 8'h9e;    Green = 8'h9e;    Blue = 8'ha6;
end 12'ha56:    begin Red = 8'hc2;    Green = 8'hbd;    Blue = 8'hc1;
end 12'ha57:    begin Red = 8'hb9;    Green = 8'hbb;    Blue = 8'hd1;
end 12'ha58:    begin Red = 8'heb;    Green = 8'hd8;    Blue = 8'hc1;
end 12'ha59:    begin Red = 8'h06;    Green = 8'hc5;    Blue = 8'h2f;
end 12'ha5a:    begin Red = 8'h05;    Green = 8'hf4;    Blue = 8'h48;
end 12'ha5b:    begin Red = 8'hfe;    Green = 8'hec;    Blue = 8'he0;
end 12'ha5c:    begin Red = 8'h73;    Green = 8'h7c;    Blue = 8'h7b;
end 12'ha5d:    begin Red = 8'haf;    Green = 8'h82;    Blue = 8'h53;
end 12'ha5e:    begin Red = 8'ha1;    Green = 8'h76;    Blue = 8'h45;
end 12'ha5f:    begin Red = 8'hf2;    Green = 8'he9;    Blue = 8'hd8;
end 12'ha60:    begin Red = 8'he2;    Green = 8'hcd;    Blue = 8'hb8;
end 12'ha61:    begin Red = 8'hc8;    Green = 8'hb3;    Blue = 8'h9e;
end 12'ha62:    begin Red = 8'h01;    Green = 8'h91;    Blue = 8'h6d;
end 12'ha63:    begin Red = 8'he0;    Green = 8'hc5;    Blue = 8'h9a;
end 12'ha64:    begin Red = 8'h76;    Green = 8'h9f;    Blue = 8'h72;
end 12'ha65:    begin Red = 8'hc8;    Green = 8'h9c;    Blue = 8'h70;
end 12'ha66:    begin Red = 8'hf1;    Green = 8'hca;    Blue = 8'h92;
end 12'ha67:    begin Red = 8'hde;    Green = 8'hbb;    Blue = 8'h82;
end 12'ha68:    begin Red = 8'hd2;    Green = 8'ha7;    Blue = 8'h71;
end 12'ha69:    begin Red = 8'hbb;    Green = 8'hb2;    Blue = 8'h9e;
end 12'ha6a:    begin Red = 8'hd1;    Green = 8'haf;    Blue = 8'h7c;
end 12'ha6b:    begin Red = 8'he1;    Green = 8'hd3;    Blue = 8'hb7;
end 12'ha6c:    begin Red = 8'hc7;    Green = 8'hd7;    Blue = 8'h9a;
end 12'ha6d:    begin Red = 8'h97;    Green = 8'h92;    Blue = 8'h6d;
end 12'ha6e:    begin Red = 8'h61;    Green = 8'h48;    Blue = 8'h3a;
end 12'ha6f:    begin Red = 8'hab;    Green = 8'h9f;    Blue = 8'h90;
end 12'ha70:    begin Red = 8'hb3;    Green = 8'h87;    Blue = 8'h6c;
end 12'ha71:    begin Red = 8'h46;    Green = 8'h43;    Blue = 8'h2a;
end 12'ha72:    begin Red = 8'hcf;    Green = 8'ha4;    Blue = 8'h76;
end 12'ha73:    begin Red = 8'h7c;    Green = 8'h63;    Blue = 8'h34;
end 12'ha74:    begin Red = 8'h73;    Green = 8'h77;    Blue = 8'h61;
end 12'ha75:    begin Red = 8'h80;    Green = 8'h87;    Blue = 8'h6f;
end 12'ha76:    begin Red = 8'hf8;    Green = 8'h99;    Blue = 8'h6b;
end 12'ha77:    begin Red = 8'h94;    Green = 8'h72;    Blue = 8'h3e;
end 12'ha78:    begin Red = 8'h92;    Green = 8'h76;    Blue = 8'h46;
end 12'ha79:    begin Red = 8'h8e;    Green = 8'h9f;    Blue = 8'h86;
end 12'ha7a:    begin Red = 8'hb4;    Green = 8'hb9;    Blue = 8'h82;
end 12'ha7b:    begin Red = 8'hc1;    Green = 8'hd5;    Blue = 8'hab;
end 12'ha7c:    begin Red = 8'hc9;    Green = 8'hb2;    Blue = 8'h84;
end 12'ha7d:    begin Red = 8'hd5;    Green = 8'h83;    Blue = 8'h49;
end 12'ha7e:    begin Red = 8'hbb;    Green = 8'hc1;    Blue = 8'h99;
end 12'ha7f:    begin Red = 8'h8b;    Green = 8'h61;    Blue = 8'h42;
end 12'ha80:    begin Red = 8'ha7;    Green = 8'h98;    Blue = 8'h8c;
end 12'ha81:    begin Red = 8'h3a;    Green = 8'h28;    Blue = 8'h1d;
end 12'ha82:    begin Red = 8'h36;    Green = 8'h23;    Blue = 8'h1c;
end 12'ha83:    begin Red = 8'hc4;    Green = 8'h64;    Blue = 8'h33;
end 12'ha84:    begin Red = 8'he5;    Green = 8'h95;    Blue = 8'h63;
end 12'ha85:    begin Red = 8'hbc;    Green = 8'hb3;    Blue = 8'h94;
end 12'ha86:    begin Red = 8'h0b;    Green = 8'h87;    Blue = 8'h4c;
end 12'ha87:    begin Red = 8'hc7;    Green = 8'h7f;    Blue = 8'h17;
end 12'ha88:    begin Red = 8'h0c;    Green = 8'ha7;    Blue = 8'hec;
end 12'ha89:    begin Red = 8'h67;    Green = 8'ha3;    Blue = 8'h5f;
end 12'ha8a:    begin Red = 8'h8a;    Green = 8'h59;    Blue = 8'h30;
end 12'ha8b:    begin Red = 8'h5e;    Green = 8'h7a;    Blue = 8'h41;
end 12'ha8c:    begin Red = 8'h64;    Green = 8'h9e;    Blue = 8'h55;
end 12'ha8d:    begin Red = 8'hd2;    Green = 8'hb6;    Blue = 8'h90;
end 12'ha8e:    begin Red = 8'hb0;    Green = 8'hb1;    Blue = 8'h91;
end 12'ha8f:    begin Red = 8'hc3;    Green = 8'hc4;    Blue = 8'ha1;
end 12'ha90:    begin Red = 8'h6c;    Green = 8'h5d;    Blue = 8'h3f;
end 12'ha91:    begin Red = 8'he6;    Green = 8'h96;    Blue = 8'h57;
end 12'ha92:    begin Red = 8'hdd;    Green = 8'h9d;    Blue = 8'h53;
end 12'ha93:    begin Red = 8'he7;    Green = 8'h98;    Blue = 8'h6a;
end 12'ha94:    begin Red = 8'hd9;    Green = 8'he2;    Blue = 8'hc6;
end 12'ha95:    begin Red = 8'hda;    Green = 8'hde;    Blue = 8'hbd;
end 12'ha96:    begin Red = 8'hdf;    Green = 8'h99;    Blue = 8'h72;
end 12'ha97:    begin Red = 8'hbc;    Green = 8'h82;    Blue = 8'h11;
end 12'ha98:    begin Red = 8'hc1;    Green = 8'h7c;    Blue = 8'h17;
end 12'ha99:    begin Red = 8'h0c;    Green = 8'h97;    Blue = 8'hce;
end 12'ha9a:    begin Red = 8'h6f;    Green = 8'ha2;    Blue = 8'h68;
end 12'ha9b:    begin Red = 8'ha2;    Green = 8'h98;    Blue = 8'h8a;
end 12'ha9c:    begin Red = 8'hb4;    Green = 8'hb0;    Blue = 8'h9e;
end 12'ha9d:    begin Red = 8'h67;    Green = 8'h64;    Blue = 8'h3c;
end 12'ha9e:    begin Red = 8'hdb;    Green = 8'h8a;    Blue = 8'h4e;
end 12'ha9f:    begin Red = 8'he3;    Green = 8'h9d;    Blue = 8'h6a;
end 12'haa0:    begin Red = 8'hed;    Green = 8'h94;    Blue = 8'h21;
end 12'haa1:    begin Red = 8'hb8;    Green = 8'h76;    Blue = 8'h1c;
end 12'haa2:    begin Red = 8'hc2;    Green = 8'h7d;    Blue = 8'h1c;
end 12'haa3:    begin Red = 8'hc9;    Green = 8'haf;    Blue = 8'h8a;
end 12'haa4:    begin Red = 8'h70;    Green = 8'h57;    Blue = 8'h32;
end 12'haa5:    begin Red = 8'h92;    Green = 8'h70;    Blue = 8'h44;
end 12'haa6:    begin Red = 8'hd4;    Green = 8'he9;    Blue = 8'hf0;
end 12'haa7:    begin Red = 8'hb3;    Green = 8'hbc;    Blue = 8'h99;
end 12'haa8:    begin Red = 8'hb5;    Green = 8'hb6;    Blue = 8'h96;
end 12'haa9:    begin Red = 8'hf1;    Green = 8'h99;    Blue = 8'h11;
end 12'haaa:    begin Red = 8'hb2;    Green = 8'h87;    Blue = 8'h58;
end 12'haab:    begin Red = 8'h37;    Green = 8'h1d;    Blue = 8'h1f;
end 12'haac:    begin Red = 8'h8a;    Green = 8'h7a;    Blue = 8'h51;
end 12'haad:    begin Red = 8'hae;    Green = 8'hb7;    Blue = 8'h8c;
end 12'haae:    begin Red = 8'haf;    Green = 8'hc3;    Blue = 8'h82;
end 12'haaf:    begin Red = 8'hef;    Green = 8'h9a;    Blue = 8'h17;
end 12'hab0:    begin Red = 8'h73;    Green = 8'h6c;    Blue = 8'h4a;
end 12'hab1:    begin Red = 8'hfa;    Green = 8'hdc;    Blue = 8'ha8;
end 12'hab2:    begin Red = 8'h00;    Green = 8'h18;    Blue = 8'h50;
end 12'hab3:    begin Red = 8'hf6;    Green = 8'hf4;    Blue = 8'hd1;
end 12'hab4:    begin Red = 8'h66;    Green = 8'h64;    Blue = 8'h45;
end 12'hab5:    begin Red = 8'ha6;    Green = 8'hac;    Blue = 8'h77;
end 12'hab6:    begin Red = 8'hce;    Green = 8'hcb;    Blue = 8'h9c;
end 12'hab7:    begin Red = 8'had;    Green = 8'ha0;    Blue = 8'h8b;
end 12'hab8:    begin Red = 8'h0e;    Green = 8'h68;    Blue = 8'h50;
end 12'hab9:    begin Red = 8'he6;    Green = 8'h90;    Blue = 8'h1d;
end 12'haba:    begin Red = 8'hdc;    Green = 8'h95;    Blue = 8'h21;
end 12'habb:    begin Red = 8'h99;    Green = 8'h8a;    Blue = 8'h7f;
end 12'habc:    begin Red = 8'h00;    Green = 8'h1b;    Blue = 8'he0;
end 12'habd:    begin Red = 8'hd7;    Green = 8'hd6;    Blue = 8'hb2;
end 12'habe:    begin Red = 8'hf5;    Green = 8'had;    Blue = 8'h70;
end 12'habf:    begin Red = 8'h7a;    Green = 8'h76;    Blue = 8'h6e;
end 12'hac0:    begin Red = 8'h6a;    Green = 8'h47;    Blue = 8'h1a;
end 12'hac1:    begin Red = 8'hff;    Green = 8'hab;    Blue = 8'h67;
end 12'hac2:    begin Red = 8'hff;    Green = 8'had;    Blue = 8'h6c;
end 12'hac3:    begin Red = 8'hff;    Green = 8'haa;    Blue = 8'h62;
end 12'hac4:    begin Red = 8'hdb;    Green = 8'hdb;    Blue = 8'hb2;
end 12'hac5:    begin Red = 8'h6c;    Green = 8'h71;    Blue = 8'h4d;
end 12'hac6:    begin Red = 8'h0e;    Green = 8'ha8;    Blue = 8'h74;
end 12'hac7:    begin Red = 8'hfd;    Green = 8'h9c;    Blue = 8'h1f;
end 12'hac8:    begin Red = 8'h0c;    Green = 8'h67;    Blue = 8'hbe;
end 12'hac9:    begin Red = 8'h97;    Green = 8'h6e;    Blue = 8'h32;
end 12'haca:    begin Red = 8'h48;    Green = 8'h4c;    Blue = 8'h37;
end 12'hacb:    begin Red = 8'h49;    Green = 8'h52;    Blue = 8'h39;
end 12'hacc:    begin Red = 8'hb4;    Green = 8'h9f;    Blue = 8'h7d;
end 12'hacd:    begin Red = 8'h61;    Green = 8'h60;    Blue = 8'h43;
end 12'hace:    begin Red = 8'hc3;    Green = 8'h6d;    Blue = 8'h2b;
end 12'hacf:    begin Red = 8'he4;    Green = 8'h93;    Blue = 8'h68;
end 12'had0:    begin Red = 8'hbd;    Green = 8'hb0;    Blue = 8'h8f;
end 12'had1:    begin Red = 8'he8;    Green = 8'h97;    Blue = 8'h21;
end 12'had2:    begin Red = 8'hfc;    Green = 8'h9e;    Blue = 8'h10;
end 12'had3:    begin Red = 8'hd3;    Green = 8'h80;    Blue = 8'h14;
end 12'had4:    begin Red = 8'h3f;    Green = 8'h4f;    Blue = 8'h2c;
end 12'had5:    begin Red = 8'h3d;    Green = 8'h4f;    Blue = 8'h3a;
end 12'had6:    begin Red = 8'h4d;    Green = 8'h5d;    Blue = 8'h3a;
end 12'had7:    begin Red = 8'h51;    Green = 8'h38;    Blue = 8'h1e;
end 12'had8:    begin Red = 8'h01;    Green = 8'hc1;    Blue = 8'h00;
end 12'had9:    begin Red = 8'hdb;    Green = 8'hc7;    Blue = 8'h96;
end 12'hada:    begin Red = 8'hf5;    Green = 8'hdb;    Blue = 8'hba;
end 12'hadb:    begin Red = 8'hbe;    Green = 8'h97;    Blue = 8'h50;
end 12'hadc:    begin Red = 8'hb9;    Green = 8'h95;    Blue = 8'h4a;
end 12'hadd:    begin Red = 8'hbc;    Green = 8'h90;    Blue = 8'h44;
end 12'hade:    begin Red = 8'h51;    Green = 8'h3d;    Blue = 8'h2b;
end 12'hadf:    begin Red = 8'hd8;    Green = 8'hbe;    Blue = 8'h97;
end 12'hae0:    begin Red = 8'h71;    Green = 8'h5f;    Blue = 8'h4b;
end 12'hae1:    begin Red = 8'h04;    Green = 8'he3;    Blue = 8'h7e;
end 12'hae2:    begin Red = 8'h03;    Green = 8'h72;    Blue = 8'h68;
end 12'hae3:    begin Red = 8'h02;    Green = 8'he1;    Blue = 8'hd9;
end 12'hae4:    begin Red = 8'h00;    Green = 8'h15;    Blue = 8'h00;
end 12'hae5:    begin Red = 8'hff;    Green = 8'hed;    Blue = 8'hd1;
end 12'hae6:    begin Red = 8'hdb;    Green = 8'hc2;    Blue = 8'h9d;
end 12'hae7:    begin Red = 8'h8d;    Green = 8'h7f;    Blue = 8'h76;
end 12'hae8:    begin Red = 8'hbb;    Green = 8'h8f;    Blue = 8'h2b;
end 12'hae9:    begin Red = 8'hb4;    Green = 8'h92;    Blue = 8'h3f;
end 12'haea:    begin Red = 8'hc3;    Green = 8'h9c;    Blue = 8'h44;
end 12'haeb:    begin Red = 8'hbe;    Green = 8'h99;    Blue = 8'h45;
end 12'haec:    begin Red = 8'hc5;    Green = 8'ha0;    Blue = 8'h4d;
end 12'haed:    begin Red = 8'hea;    Green = 8'h93;    Blue = 8'h51;
end 12'haee:    begin Red = 8'hd3;    Green = 8'he5;    Blue = 8'hc2;
end 12'haef:    begin Red = 8'hd7;    Green = 8'he3;    Blue = 8'hcc;
end 12'haf0:    begin Red = 8'hf1;    Green = 8'hdb;    Blue = 8'hb4;
end 12'haf1:    begin Red = 8'hff;    Green = 8'hd2;    Blue = 8'h9a;
end 12'haf2:    begin Red = 8'he7;    Green = 8'hc3;    Blue = 8'h9a;
end 12'haf3:    begin Red = 8'h9d;    Green = 8'h7f;    Blue = 8'h3c;
end 12'haf4:    begin Red = 8'h96;    Green = 8'h77;    Blue = 8'h36;
end 12'haf5:    begin Red = 8'had;    Green = 8'hb9;    Blue = 8'h9c;
end 12'haf6:    begin Red = 8'h58;    Green = 8'h40;    Blue = 8'h1e;
end 12'haf7:    begin Red = 8'h94;    Green = 8'h80;    Blue = 8'h6c;
end 12'haf8:    begin Red = 8'h03;    Green = 8'h12;    Blue = 8'h68;
end 12'haf9:    begin Red = 8'h31;    Green = 8'h34;    Blue = 8'h32;
end 12'hafa:    begin Red = 8'h5b;    Green = 8'h3c;    Blue = 8'h18;
end 12'hafb:    begin Red = 8'h47;    Green = 8'h32;    Blue = 8'h3c;
end 12'hafc:    begin Red = 8'h00;    Green = 8'h1b;    Blue = 8'h70;
end 12'hafd:    begin Red = 8'hec;    Green = 8'hbd;    Blue = 8'h83;
end 12'hafe:    begin Red = 8'h42;    Green = 8'h36;    Blue = 8'h31;
end 12'haff:    begin Red = 8'h30;    Green = 8'h2a;    Blue = 8'h2b;
end 12'hb00:    begin Red = 8'h8d;    Green = 8'h77;    Blue = 8'h62;
end 12'hb01:    begin Red = 8'h02;    Green = 8'h91;    Blue = 8'h79;
end 12'hb02:    begin Red = 8'hb4;    Green = 8'h8f;    Blue = 8'h58;
end 12'hb03:    begin Red = 8'he5;    Green = 8'hf5;    Blue = 8'hd3;
end 12'hb04:    begin Red = 8'heb;    Green = 8'hef;    Blue = 8'hca;
end 12'hb05:    begin Red = 8'hed;    Green = 8'hf0;    Blue = 8'hdf;
end 12'hb06:    begin Red = 8'h81;    Green = 8'h72;    Blue = 8'h63;
end 12'hb07:    begin Red = 8'h7b;    Green = 8'h6f;    Blue = 8'h6a;
end 12'hb08:    begin Red = 8'h82;    Green = 8'h58;    Blue = 8'h2a;
end 12'hb09:    begin Red = 8'h6f;    Green = 8'h49;    Blue = 8'h12;
end 12'hb0a:    begin Red = 8'hf7;    Green = 8'he9;    Blue = 8'hc5;
end 12'hb0b:    begin Red = 8'hc4;    Green = 8'hc1;    Blue = 8'ha9;
end 12'hb0c:    begin Red = 8'h63;    Green = 8'h5a;    Blue = 8'h56;
end 12'hb0d:    begin Red = 8'hb4;    Green = 8'h92;    Blue = 8'h45;
end 12'hb0e:    begin Red = 8'h9b;    Green = 8'h4d;    Blue = 8'h2e;
end 12'hb0f:    begin Red = 8'h91;    Green = 8'h4f;    Blue = 8'h2e;
end 12'hb10:    begin Red = 8'h91;    Green = 8'h57;    Blue = 8'h2a;
end 12'hb11:    begin Red = 8'h01;    Green = 8'h21;    Blue = 8'h00;
end 12'hb12:    begin Red = 8'haf;    Green = 8'h78;    Blue = 8'h4a;
end 12'hb13:    begin Red = 8'hb2;    Green = 8'h68;    Blue = 8'h3e;
end 12'hb14:    begin Red = 8'hb8;    Green = 8'hbe;    Blue = 8'h88;
end 12'hb15:    begin Red = 8'hfe;    Green = 8'hf5;    Blue = 8'hd1;
end 12'hb16:    begin Red = 8'hd8;    Green = 8'hde;    Blue = 8'hab;
end 12'hb17:    begin Red = 8'hbd;    Green = 8'h9c;    Blue = 8'h6e;
end 12'hb18:    begin Red = 8'h69;    Green = 8'h56;    Blue = 8'h2f;
end 12'hb19:    begin Red = 8'hc9;    Green = 8'hb9;    Blue = 8'h93;
end 12'hb1a:    begin Red = 8'h4d;    Green = 8'h49;    Blue = 8'h43;
end 12'hb1b:    begin Red = 8'hcd;    Green = 8'hb8;    Blue = 8'h8a;
end 12'hb1c:    begin Red = 8'h4e;    Green = 8'h40;    Blue = 8'h36;
end 12'hb1d:    begin Red = 8'ha7;    Green = 8'h8b;    Blue = 8'h78;
end 12'hb1e:    begin Red = 8'h86;    Green = 8'h72;    Blue = 8'h62;
end 12'hb1f:    begin Red = 8'hbc;    Green = 8'h94;    Blue = 8'h2f;
end 12'hb20:    begin Red = 8'h94;    Green = 8'h6f;    Blue = 8'h25;
end 12'hb21:    begin Red = 8'hca;    Green = 8'ha0;    Blue = 8'h4a;
end 12'hb22:    begin Red = 8'hd0;    Green = 8'ha9;    Blue = 8'h58;
end 12'hb23:    begin Red = 8'h87;    Green = 8'h6b;    Blue = 8'h26;
end 12'hb24:    begin Red = 8'h96;    Green = 8'h46;    Blue = 8'h27;
end 12'hb25:    begin Red = 8'ha4;    Green = 8'h5c;    Blue = 8'h2d;
end 12'hb26:    begin Red = 8'hdb;    Green = 8'h8b;    Blue = 8'h5c;
end 12'hb27:    begin Red = 8'h66;    Green = 8'h5e;    Blue = 8'h41;
end 12'hb28:    begin Red = 8'hba;    Green = 8'h70;    Blue = 8'h42;
end 12'hb29:    begin Red = 8'hc1;    Green = 8'h76;    Blue = 8'h36;
end 12'hb2a:    begin Red = 8'hfe;    Green = 8'hef;    Blue = 8'hbb;
end 12'hb2b:    begin Red = 8'h76;    Green = 8'h79;    Blue = 8'h54;
end 12'hb2c:    begin Red = 8'h47;    Green = 8'h33;    Blue = 8'h22;
end 12'hb2d:    begin Red = 8'h03;    Green = 8'he2;    Blue = 8'hde;
end 12'hb2e:    begin Red = 8'h73;    Green = 8'h5b;    Blue = 8'h27;
end 12'hb2f:    begin Red = 8'h6e;    Green = 8'h53;    Blue = 8'h45;
end 12'hb30:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'h3f;
end 12'hb31:    begin Red = 8'h93;    Green = 8'h84;    Blue = 8'h67;
end 12'hb32:    begin Red = 8'h54;    Green = 8'h48;    Blue = 8'h2a;
end 12'hb33:    begin Red = 8'h81;    Green = 8'h65;    Blue = 8'h52;
end 12'hb34:    begin Red = 8'h66;    Green = 8'h4c;    Blue = 8'h44;
end 12'hb35:    begin Red = 8'hb1;    Green = 8'h8c;    Blue = 8'h3b;
end 12'hb36:    begin Red = 8'hc2;    Green = 8'h8f;    Blue = 8'h40;
end 12'hb37:    begin Red = 8'hc3;    Green = 8'hb6;    Blue = 8'h93;
end 12'hb38:    begin Red = 8'h00;    Green = 8'h0f;    Blue = 8'h04;
end 12'hb39:    begin Red = 8'h00;    Green = 8'h17;    Blue = 8'h96;
end 12'hb3a:    begin Red = 8'h00;    Green = 8'h03;    Blue = 8'h00;
end 12'hb3b:    begin Red = 8'h65;    Green = 8'h4a;    Blue = 8'h2e;
end 12'hb3c:    begin Red = 8'hb0;    Green = 8'h86;    Blue = 8'h2b;
end 12'hb3d:    begin Red = 8'ha3;    Green = 8'h80;    Blue = 8'h37;
end 12'hb3e:    begin Red = 8'hb5;    Green = 8'h85;    Blue = 8'h34;
end 12'hb3f:    begin Red = 8'hbb;    Green = 8'ha8;    Blue = 8'h70;
end 12'hb40:    begin Red = 8'h65;    Green = 8'h61;    Blue = 8'h4e;
end 12'hb41:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'h9d;
end 12'hb42:    begin Red = 8'h33;    Green = 8'h24;    Blue = 8'h10;
end 12'hb43:    begin Red = 8'h00;    Green = 8'h0f;    Blue = 8'hf3;
end 12'hb44:    begin Red = 8'hbf;    Green = 8'hb2;    Blue = 8'h81;
end 12'hb45:    begin Red = 8'ha3;    Green = 8'h9a;    Blue = 8'h6a;
end 12'hb46:    begin Red = 8'h92;    Green = 8'h8c;    Blue = 8'h65;
end 12'hb47:    begin Red = 8'h62;    Green = 8'h4c;    Blue = 8'h4f;
end 12'hb48:    begin Red = 8'h56;    Green = 8'h54;    Blue = 8'h3f;
end 12'hb49:    begin Red = 8'h8e;    Green = 8'h6e;    Blue = 8'h1c;
end 12'hb4a:    begin Red = 8'ha5;    Green = 8'h86;    Blue = 8'h3f;
end 12'hb4b:    begin Red = 8'h9d;    Green = 8'h7e;    Blue = 8'h34;
end 12'hb4c:    begin Red = 8'hc0;    Green = 8'h8d;    Blue = 8'h51;
end 12'hb4d:    begin Red = 8'hc5;    Green = 8'h96;    Blue = 8'h5a;
end 12'hb4e:    begin Red = 8'had;    Green = 8'h7d;    Blue = 8'h48;
end 12'hb4f:    begin Red = 8'hb3;    Green = 8'h87;    Blue = 8'h42;
end 12'hb50:    begin Red = 8'hb7;    Green = 8'h8e;    Blue = 8'h52;
end 12'hb51:    begin Red = 8'hb2;    Green = 8'h87;    Blue = 8'h47;
end 12'hb52:    begin Red = 8'hb7;    Green = 8'h8c;    Blue = 8'h4d;
end 12'hb53:    begin Red = 8'h81;    Green = 8'h5e;    Blue = 8'h37;
end 12'hb54:    begin Red = 8'h5d;    Green = 8'h49;    Blue = 8'h4d;
end 12'hb55:    begin Red = 8'h58;    Green = 8'h4e;    Blue = 8'h48;
end 12'hb56:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h95;
end 12'hb57:    begin Red = 8'h04;    Green = 8'hf2;    Blue = 8'he6;
end 12'hb58:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'hff;
end 12'hb59:    begin Red = 8'h53;    Green = 8'h39;    Blue = 8'h31;
end 12'hb5a:    begin Red = 8'h82;    Green = 8'h57;    Blue = 8'h48;
end 12'hb5b:    begin Red = 8'h82;    Green = 8'h5c;    Blue = 8'h48;
end 12'hb5c:    begin Red = 8'h86;    Green = 8'h67;    Blue = 8'h21;
end 12'hb5d:    begin Red = 8'hae;    Green = 8'h87;    Blue = 8'h3b;
end 12'hb5e:    begin Red = 8'hb0;    Green = 8'h86;    Blue = 8'h35;
end 12'hb5f:    begin Red = 8'had;    Green = 8'h87;    Blue = 8'h40;
end 12'hb60:    begin Red = 8'h04;    Green = 8'h53;    Blue = 8'h18;
end 12'hb61:    begin Red = 8'h04;    Green = 8'h83;    Blue = 8'h00;
end 12'hb62:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'hb6;
end 12'hb63:    begin Red = 8'h00;    Green = 8'h18;    Blue = 8'hdb;
end 12'hb64:    begin Red = 8'h3f;    Green = 8'h30;    Blue = 8'h2e;
end 12'hb65:    begin Red = 8'h53;    Green = 8'h41;    Blue = 8'h36;
end 12'hb66:    begin Red = 8'h02;    Green = 8'hc1;    Blue = 8'hbb;
end 12'hb67:    begin Red = 8'h6a;    Green = 8'h81;    Blue = 8'h9e;
end 12'hb68:    begin Red = 8'h6f;    Green = 8'h83;    Blue = 8'hb5;
end 12'hb69:    begin Red = 8'h94;    Green = 8'h6d;    Blue = 8'h2b;
end 12'hb6a:    begin Red = 8'h6e;    Green = 8'h93;    Blue = 8'hc9;
end 12'hb6b:    begin Red = 8'h6e;    Green = 8'h82;    Blue = 8'ha8;
end 12'hb6c:    begin Red = 8'h77;    Green = 8'h91;    Blue = 8'hcb;
end 12'hb6d:    begin Red = 8'h00;    Green = 8'h0c;    Blue = 8'h7b;
end 12'hb6e:    begin Red = 8'hd7;    Green = 8'ha9;    Blue = 8'h6a;
end 12'hb6f:    begin Red = 8'hee;    Green = 8'hc3;    Blue = 8'h7f;
end 12'hb70:    begin Red = 8'he9;    Green = 8'hc0;    Blue = 8'h7b;
end 12'hb71:    begin Red = 8'hdf;    Green = 8'he0;    Blue = 8'hc6;
end 12'hb72:    begin Red = 8'he2;    Green = 8'hb9;    Blue = 8'h76;
end 12'hb73:    begin Red = 8'hde;    Green = 8'hb3;    Blue = 8'h71;
end 12'hb74:    begin Red = 8'hb3;    Green = 8'h95;    Blue = 8'h55;
end 12'hb75:    begin Red = 8'heb;    Green = 8'hc5;    Blue = 8'h8e;
end 12'hb76:    begin Red = 8'h06;    Green = 8'h93;    Blue = 8'hb0;
end 12'hb77:    begin Red = 8'h07;    Green = 8'hf4;    Blue = 8'hf8;
end 12'hb78:    begin Red = 8'h06;    Green = 8'h94;    Blue = 8'h03;
end 12'hb79:    begin Red = 8'hca;    Green = 8'h9d;    Blue = 8'h64;
end 12'hb7a:    begin Red = 8'hd0;    Green = 8'ha6;    Blue = 8'h5f;
end 12'hb7b:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'hb8;
end 12'hb7c:    begin Red = 8'h07;    Green = 8'h94;    Blue = 8'hb9;
end 12'hb7d:    begin Red = 8'h07;    Green = 8'h44;    Blue = 8'hdd;
end 12'hb7e:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'hb5;
end 12'hb7f:    begin Red = 8'h05;    Green = 8'h22;    Blue = 8'h42;
end 12'hb80:    begin Red = 8'hbd;    Green = 8'h94;    Blue = 8'h5c;
end 12'hb81:    begin Red = 8'haf;    Green = 8'h8a;    Blue = 8'h51;
end 12'hb82:    begin Red = 8'hd4;    Green = 8'hdc;    Blue = 8'hb6;
end 12'hb83:    begin Red = 8'haa;    Green = 8'h85;    Blue = 8'h51;
end 12'hb84:    begin Red = 8'h06;    Green = 8'h23;    Blue = 8'he7;
end 12'hb85:    begin Red = 8'h05;    Green = 8'he3;    Blue = 8'hc8;
end 12'hb86:    begin Red = 8'h05;    Green = 8'hd3;    Blue = 8'he3;
end 12'hb87:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'hf5;
end 12'hb88:    begin Red = 8'hac;    Green = 8'h82;    Blue = 8'h26;
end 12'hb89:    begin Red = 8'ha8;    Green = 8'h80;    Blue = 8'h3c;
end 12'hb8a:    begin Red = 8'hd6;    Green = 8'ha7;    Blue = 8'h64;
end 12'hb8b:    begin Red = 8'h08;    Green = 8'h05;    Blue = 8'h0d;
end 12'hb8c:    begin Red = 8'h08;    Green = 8'h44;    Blue = 8'hf5;
end 12'hb8d:    begin Red = 8'h08;    Green = 8'h24;    Blue = 8'hee;
end 12'hb8e:    begin Red = 8'h06;    Green = 8'h64;    Blue = 8'h0a;
end 12'hb8f:    begin Red = 8'hcf;    Green = 8'ha7;    Blue = 8'h64;
end 12'hb90:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'h70;
end 12'hb91:    begin Red = 8'h07;    Green = 8'hb5;    Blue = 8'h07;
end 12'hb92:    begin Red = 8'h07;    Green = 8'h64;    Blue = 8'hd9;
end 12'hb93:    begin Red = 8'h07;    Green = 8'h84;    Blue = 8'hf8;
end 12'hb94:    begin Red = 8'h06;    Green = 8'h44;    Blue = 8'h2d;
end 12'hb95:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'hc7;
end 12'hb96:    begin Red = 8'h04;    Green = 8'hd2;    Blue = 8'hd2;
end 12'hb97:    begin Red = 8'h8f;    Green = 8'h6f;    Blue = 8'h69;
end 12'hb98:    begin Red = 8'h8d;    Green = 8'h6a;    Blue = 8'h66;
end 12'hb99:    begin Red = 8'h73;    Green = 8'h58;    Blue = 8'h55;
end 12'hb9a:    begin Red = 8'h8e;    Green = 8'h6a;    Blue = 8'h6d;
end 12'hb9b:    begin Red = 8'h8a;    Green = 8'h68;    Blue = 8'h61;
end 12'hb9c:    begin Red = 8'h58;    Green = 8'h3d;    Blue = 8'h48;
end 12'hb9d:    begin Red = 8'h7a;    Green = 8'h56;    Blue = 8'h5a;
end 12'hb9e:    begin Red = 8'h97;    Green = 8'h6e;    Blue = 8'h6c;
end 12'hb9f:    begin Red = 8'h8e;    Green = 8'h60;    Blue = 8'h61;
end 12'hba0:    begin Red = 8'h78;    Green = 8'h5b;    Blue = 8'h58;
end 12'hba1:    begin Red = 8'h5f;    Green = 8'h40;    Blue = 8'h4a;
end 12'hba2:    begin Red = 8'h01;    Green = 8'hc1;    Blue = 8'h5d;
end 12'hba3:    begin Red = 8'hf8;    Green = 8'heb;    Blue = 8'hcc;
end 12'hba4:    begin Red = 8'hee;    Green = 8'hc2;    Blue = 8'h85;
end 12'hba5:    begin Red = 8'h8b;    Green = 8'h55;    Blue = 8'h13;
end 12'hba6:    begin Red = 8'h06;    Green = 8'hc4;    Blue = 8'h44;
end 12'hba7:    begin Red = 8'hf6;    Green = 8'hd2;    Blue = 8'h92;
end 12'hba8:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'h98;
end 12'hba9:    begin Red = 8'h9d;    Green = 8'h7c;    Blue = 8'h49;
end 12'hbaa:    begin Red = 8'h98;    Green = 8'h6b;    Blue = 8'h3d;
end 12'hbab:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'he5;
end 12'hbac:    begin Red = 8'h78;    Green = 8'h5e;    Blue = 8'h5f;
end 12'hbad:    begin Red = 8'ha5;    Green = 8'h7c;    Blue = 8'h7a;
end 12'hbae:    begin Red = 8'ha9;    Green = 8'h85;    Blue = 8'h80;
end 12'hbaf:    begin Red = 8'ha8;    Green = 8'h7f;    Blue = 8'h72;
end 12'hbb0:    begin Red = 8'h6d;    Green = 8'h51;    Blue = 8'h58;
end 12'hbb1:    begin Red = 8'h85;    Green = 8'h68;    Blue = 8'h64;
end 12'hbb2:    begin Red = 8'h73;    Green = 8'h50;    Blue = 8'h5f;
end 12'hbb3:    begin Red = 8'h78;    Green = 8'h59;    Blue = 8'h61;
end 12'hbb4:    begin Red = 8'hb1;    Green = 8'h86;    Blue = 8'h83;
end 12'hbb5:    begin Red = 8'hac;    Green = 8'h7c;    Blue = 8'h7f;
end 12'hbb6:    begin Red = 8'hb6;    Green = 8'h89;    Blue = 8'h24;
end 12'hbb7:    begin Red = 8'h01;    Green = 8'he1;    Blue = 8'h3d;
end 12'hbb8:    begin Red = 8'hd2;    Green = 8'hc9;    Blue = 8'hab;
end 12'hbb9:    begin Red = 8'hd2;    Green = 8'hc4;    Blue = 8'ha6;
end 12'hbba:    begin Red = 8'h07;    Green = 8'hd4;    Blue = 8'hba;
end 12'hbbb:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'hf5;
end 12'hbbc:    begin Red = 8'h98;    Green = 8'h70;    Blue = 8'h38;
end 12'hbbd:    begin Red = 8'hdb;    Green = 8'hae;    Blue = 8'h68;
end 12'hbbe:    begin Red = 8'he4;    Green = 8'hba;    Blue = 8'h7b;
end 12'hbbf:    begin Red = 8'h07;    Green = 8'ha4;    Blue = 8'ha7;
end 12'hbc0:    begin Red = 8'h05;    Green = 8'hc3;    Blue = 8'h83;
end 12'hbc1:    begin Red = 8'hc8;    Green = 8'h97;    Blue = 8'h67;
end 12'hbc2:    begin Red = 8'h83;    Green = 8'h62;    Blue = 8'h32;
end 12'hbc3:    begin Red = 8'ha5;    Green = 8'h83;    Blue = 8'h4b;
end 12'hbc4:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'ha6;
end 12'hbc5:    begin Red = 8'h82;    Green = 8'h63;    Blue = 8'h5f;
end 12'hbc6:    begin Red = 8'h9f;    Green = 8'h7b;    Blue = 8'h76;
end 12'hbc7:    begin Red = 8'h73;    Green = 8'h49;    Blue = 8'h57;
end 12'hbc8:    begin Red = 8'haa;    Green = 8'h7d;    Blue = 8'h79;
end 12'hbc9:    begin Red = 8'h73;    Green = 8'h4f;    Blue = 8'h54;
end 12'hbca:    begin Red = 8'hfe;    Green = 8'hee;    Blue = 8'hb6;
end 12'hbcb:    begin Red = 8'haa;    Green = 8'h75;    Blue = 8'h7e;
end 12'hbcc:    begin Red = 8'hf7;    Green = 8'hd2;    Blue = 8'hb0;
end 12'hbcd:    begin Red = 8'h8d;    Green = 8'h6f;    Blue = 8'h2c;
end 12'hbce:    begin Red = 8'h99;    Green = 8'h74;    Blue = 8'h2a;
end 12'hbcf:    begin Red = 8'hb8;    Green = 8'h97;    Blue = 8'h45;
end 12'hbd0:    begin Red = 8'hce;    Green = 8'hcc;    Blue = 8'hb0;
end 12'hbd1:    begin Red = 8'h22;    Green = 8'h14;    Blue = 8'h12;
end 12'hbd2:    begin Red = 8'hbb;    Green = 8'hbb;    Blue = 8'ha1;
end 12'hbd3:    begin Red = 8'h08;    Green = 8'h14;    Blue = 8'hdd;
end 12'hbd4:    begin Red = 8'h08;    Green = 8'h45;    Blue = 8'h1d;
end 12'hbd5:    begin Red = 8'he4;    Green = 8'hc0;    Blue = 8'h7e;
end 12'hbd6:    begin Red = 8'hfb;    Green = 8'hd1;    Blue = 8'h91;
end 12'hbd7:    begin Red = 8'h05;    Green = 8'hc3;    Blue = 8'ha6;
end 12'hbd8:    begin Red = 8'hc8;    Green = 8'ha2;    Blue = 8'h70;
end 12'hbd9:    begin Red = 8'h05;    Green = 8'h12;    Blue = 8'hf5;
end 12'hbda:    begin Red = 8'h03;    Green = 8'hf1;    Blue = 8'hc0;
end 12'hbdb:    begin Red = 8'ha8;    Green = 8'h74;    Blue = 8'h78;
end 12'hbdc:    begin Red = 8'h22;    Green = 8'h26;    Blue = 8'h63;
end 12'hbdd:    begin Red = 8'h49;    Green = 8'h46;    Blue = 8'h75;
end 12'hbde:    begin Red = 8'h3f;    Green = 8'h46;    Blue = 8'h68;
end 12'hbdf:    begin Red = 8'h43;    Green = 8'h3d;    Blue = 8'h7c;
end 12'hbe0:    begin Red = 8'h46;    Green = 8'h4a;    Blue = 8'h6d;
end 12'hbe1:    begin Red = 8'h45;    Green = 8'h47;    Blue = 8'h67;
end 12'hbe2:    begin Red = 8'hea;    Green = 8'hdf;    Blue = 8'hbb;
end 12'hbe3:    begin Red = 8'hde;    Green = 8'hdb;    Blue = 8'hc4;
end 12'hbe4:    begin Red = 8'hcf;    Green = 8'ha9;    Blue = 8'h69;
end 12'hbe5:    begin Red = 8'hc4;    Green = 8'h9d;    Blue = 8'h64;
end 12'hbe6:    begin Red = 8'ha0;    Green = 8'h76;    Blue = 8'h77;
end 12'hbe7:    begin Red = 8'ha5;    Green = 8'h80;    Blue = 8'h7f;
end 12'hbe8:    begin Red = 8'h6c;    Green = 8'h48;    Blue = 8'h4a;
end 12'hbe9:    begin Red = 8'hff;    Green = 8'hef;    Blue = 8'haf;
end 12'hbea:    begin Red = 8'h84;    Green = 8'h63;    Blue = 8'h64;
end 12'hbeb:    begin Red = 8'h00;    Green = 8'h1a;    Blue = 8'h69;
end 12'hbec:    begin Red = 8'h25;    Green = 8'h2b;    Blue = 8'h65;
end 12'hbed:    begin Red = 8'h1e;    Green = 8'h29;    Blue = 8'h5e;
end 12'hbee:    begin Red = 8'h1b;    Green = 8'h23;    Blue = 8'h70;
end 12'hbef:    begin Red = 8'h92;    Green = 8'h8b;    Blue = 8'h85;
end 12'hbf0:    begin Red = 8'hcd;    Green = 8'hc1;    Blue = 8'ha4;
end 12'hbf1:    begin Red = 8'h2c;    Green = 8'h32;    Blue = 8'h66;
end 12'hbf2:    begin Red = 8'h29;    Green = 8'h30;    Blue = 8'h5d;
end 12'hbf3:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'h20;
end 12'hbf4:    begin Red = 8'h06;    Green = 8'h93;    Blue = 8'h62;
end 12'hbf5:    begin Red = 8'hef;    Green = 8'hc8;    Blue = 8'h80;
end 12'hbf6:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'h37;
end 12'hbf7:    begin Red = 8'hd7;    Green = 8'hb1;    Blue = 8'h71;
end 12'hbf8:    begin Red = 8'hd2;    Green = 8'hae;    Blue = 8'h6c;
end 12'hbf9:    begin Red = 8'hbb;    Green = 8'h98;    Blue = 8'h61;
end 12'hbfa:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'h93;
end 12'hbfb:    begin Red = 8'h03;    Green = 8'hc1;    Blue = 8'hd1;
end 12'hbfc:    begin Red = 8'h00;    Green = 8'h31;    Blue = 8'hf0;
end 12'hbfd:    begin Red = 8'h9b;    Green = 8'h73;    Blue = 8'h71;
end 12'hbfe:    begin Red = 8'h6f;    Green = 8'h44;    Blue = 8'h56;
end 12'hbff:    begin Red = 8'h6d;    Green = 8'h50;    Blue = 8'h4a;
end 12'hc00:    begin Red = 8'h82;    Green = 8'h5b;    Blue = 8'h64;
end 12'hc01:    begin Red = 8'ha3;    Green = 8'h7a;    Blue = 8'h6f;
end 12'hc02:    begin Red = 8'hc5;    Green = 8'hc7;    Blue = 8'ha8;
end 12'hc03:    begin Red = 8'hd1;    Green = 8'hb3;    Blue = 8'h72;
end 12'hc04:    begin Red = 8'h92;    Green = 8'h88;    Blue = 8'h7b;
end 12'hc05:    begin Red = 8'haa;    Green = 8'h7f;    Blue = 8'h34;
end 12'hc06:    begin Red = 8'ha3;    Green = 8'h87;    Blue = 8'h39;
end 12'hc07:    begin Red = 8'h9f;    Green = 8'h80;    Blue = 8'h41;
end 12'hc08:    begin Red = 8'hb9;    Green = 8'ha5;    Blue = 8'h9e;
end 12'hc09:    begin Red = 8'hb5;    Green = 8'ha7;    Blue = 8'h8c;
end 12'hc0a:    begin Red = 8'hf3;    Green = 8'hc5;    Blue = 8'h85;
end 12'hc0b:    begin Red = 8'heb;    Green = 8'hbb;    Blue = 8'h7b;
end 12'hc0c:    begin Red = 8'hde;    Green = 8'hb3;    Blue = 8'h79;
end 12'hc0d:    begin Red = 8'ha2;    Green = 8'h7d;    Blue = 8'h48;
end 12'hc0e:    begin Red = 8'hb0;    Green = 8'h8c;    Blue = 8'h5d;
end 12'hc0f:    begin Red = 8'hf9;    Green = 8'hfc;    Blue = 8'hca;
end 12'hc10:    begin Red = 8'hf7;    Green = 8'he8;    Blue = 8'hbc;
end 12'hc11:    begin Red = 8'hed;    Green = 8'he5;    Blue = 8'ha8;
end 12'hc12:    begin Red = 8'hfc;    Green = 8'hfc;    Blue = 8'hd2;
end 12'hc13:    begin Red = 8'h52;    Green = 8'h52;    Blue = 8'h52;
end 12'hc14:    begin Red = 8'h64;    Green = 8'h67;    Blue = 8'h64;
end 12'hc15:    begin Red = 8'h7b;    Green = 8'h4e;    Blue = 8'h7c;
end 12'hc16:    begin Red = 8'hcd;    Green = 8'ha4;    Blue = 8'h3b;
end 12'hc17:    begin Red = 8'h65;    Green = 8'h60;    Blue = 8'h55;
end 12'hc18:    begin Red = 8'hd8;    Green = 8'haf;    Blue = 8'h61;
end 12'hc19:    begin Red = 8'he3;    Green = 8'hb4;    Blue = 8'h77;
end 12'hc1a:    begin Red = 8'h4e;    Green = 8'h32;    Blue = 8'h29;
end 12'hc1b:    begin Red = 8'hd4;    Green = 8'he1;    Blue = 8'hb7;
end 12'hc1c:    begin Red = 8'h80;    Green = 8'h8c;    Blue = 8'h70;
end 12'hc1d:    begin Red = 8'hab;    Green = 8'h8b;    Blue = 8'h4c;
end 12'hc1e:    begin Red = 8'hd4;    Green = 8'hc6;    Blue = 8'h9d;
end 12'hc1f:    begin Red = 8'h7c;    Green = 8'h74;    Blue = 8'h67;
end 12'hc20:    begin Red = 8'h97;    Green = 8'h8e;    Blue = 8'h85;
end 12'hc21:    begin Red = 8'h7f;    Green = 8'h59;    Blue = 8'h77;
end 12'hc22:    begin Red = 8'h80;    Green = 8'h50;    Blue = 8'h6d;
end 12'hc23:    begin Red = 8'hc7;    Green = 8'h9d;    Blue = 8'h3d;
end 12'hc24:    begin Red = 8'hc1;    Green = 8'h98;    Blue = 8'h4a;
end 12'hc25:    begin Red = 8'h00;    Green = 8'h10;    Blue = 8'h48;
end 12'hc26:    begin Red = 8'h01;    Green = 8'ha1;    Blue = 8'h5e;
end 12'hc27:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'h93;
end 12'hc28:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'h50;
end 12'hc29:    begin Red = 8'hd5;    Green = 8'hce;    Blue = 8'hac;
end 12'hc2a:    begin Red = 8'he8;    Green = 8'hb9;    Blue = 8'h76;
end 12'hc2b:    begin Red = 8'hca;    Green = 8'h9c;    Blue = 8'h5a;
end 12'hc2c:    begin Red = 8'hd4;    Green = 8'hdf;    Blue = 8'hb0;
end 12'hc2d:    begin Red = 8'h96;    Green = 8'h66;    Blue = 8'h86;
end 12'hc2e:    begin Red = 8'h80;    Green = 8'h52;    Blue = 8'h76;
end 12'hc2f:    begin Red = 8'h81;    Green = 8'h47;    Blue = 8'h7b;
end 12'hc30:    begin Red = 8'hbb;    Green = 8'h8d;    Blue = 8'h34;
end 12'hc31:    begin Red = 8'ha4;    Green = 8'h83;    Blue = 8'h2f;
end 12'hc32:    begin Red = 8'h20;    Green = 8'h20;    Blue = 8'h15;
end 12'hc33:    begin Red = 8'hf3;    Green = 8'hcb;    Blue = 8'h89;
end 12'hc34:    begin Red = 8'he1;    Green = 8'hc4;    Blue = 8'h8a;
end 12'hc35:    begin Red = 8'ha0;    Green = 8'h91;    Blue = 8'h4c;
end 12'hc36:    begin Red = 8'ha3;    Green = 8'h8c;    Blue = 8'h4a;
end 12'hc37:    begin Red = 8'hc3;    Green = 8'ha6;    Blue = 8'h60;
end 12'hc38:    begin Red = 8'hbc;    Green = 8'ha2;    Blue = 8'h57;
end 12'hc39:    begin Red = 8'hbf;    Green = 8'h9e;    Blue = 8'h5d;
end 12'hc3a:    begin Red = 8'hc8;    Green = 8'ha9;    Blue = 8'h62;
end 12'hc3b:    begin Red = 8'hc6;    Green = 8'hae;    Blue = 8'h64;
end 12'hc3c:    begin Red = 8'hc6;    Green = 8'ha7;    Blue = 8'h6b;
end 12'hc3d:    begin Red = 8'ha0;    Green = 8'h87;    Blue = 8'h48;
end 12'hc3e:    begin Red = 8'hb7;    Green = 8'ha1;    Blue = 8'h59;
end 12'hc3f:    begin Red = 8'hbe;    Green = 8'ha4;    Blue = 8'h5d;
end 12'hc40:    begin Red = 8'hbd;    Green = 8'hab;    Blue = 8'h5f;
end 12'hc41:    begin Red = 8'hc0;    Green = 8'ha7;    Blue = 8'h56;
end 12'hc42:    begin Red = 8'ha1;    Green = 8'h9d;    Blue = 8'h8e;
end 12'hc43:    begin Red = 8'h9e;    Green = 8'h8d;    Blue = 8'h87;
end 12'hc44:    begin Red = 8'haf;    Green = 8'hb7;    Blue = 8'hb2;
end 12'hc45:    begin Red = 8'hdf;    Green = 8'he9;    Blue = 8'hd3;
end 12'hc46:    begin Red = 8'hda;    Green = 8'he4;    Blue = 8'hb6;
end 12'hc47:    begin Red = 8'h9e;    Green = 8'h73;    Blue = 8'h93;
end 12'hc48:    begin Red = 8'ha6;    Green = 8'h77;    Blue = 8'h97;
end 12'hc49:    begin Red = 8'ha4;    Green = 8'h71;    Blue = 8'h92;
end 12'hc4a:    begin Red = 8'h78;    Green = 8'h52;    Blue = 8'h71;
end 12'hc4b:    begin Red = 8'h9e;    Green = 8'h67;    Blue = 8'h83;
end 12'hc4c:    begin Red = 8'hbf;    Green = 8'h81;    Blue = 8'hb7;
end 12'hc4d:    begin Red = 8'h97;    Green = 8'h6d;    Blue = 8'h91;
end 12'hc4e:    begin Red = 8'h92;    Green = 8'h5f;    Blue = 8'h81;
end 12'hc4f:    begin Red = 8'h8c;    Green = 8'h4f;    Blue = 8'h8b;
end 12'hc50:    begin Red = 8'h81;    Green = 8'h54;    Blue = 8'h68;
end 12'hc51:    begin Red = 8'h85;    Green = 8'h56;    Blue = 8'h6d;
end 12'hc52:    begin Red = 8'h8e;    Green = 8'h6d;    Blue = 8'h24;
end 12'hc53:    begin Red = 8'h0c;    Green = 8'he7;    Blue = 8'h40;
end 12'hc54:    begin Red = 8'hcd;    Green = 8'h79;    Blue = 8'h13;
end 12'hc55:    begin Red = 8'h0c;    Green = 8'ha7;    Blue = 8'h8f;
end 12'hc56:    begin Red = 8'h0c;    Green = 8'h27;    Blue = 8'h00;
end 12'hc57:    begin Red = 8'ha5;    Green = 8'h84;    Blue = 8'h46;
end 12'hc58:    begin Red = 8'hfa;    Green = 8'he4;    Blue = 8'h9e;
end 12'hc59:    begin Red = 8'hbe;    Green = 8'h86;    Blue = 8'ha9;
end 12'hc5a:    begin Red = 8'h85;    Green = 8'h4c;    Blue = 8'h85;
end 12'hc5b:    begin Red = 8'ha5;    Green = 8'ha6;    Blue = 8'h79;
end 12'hc5c:    begin Red = 8'h0b;    Green = 8'hf7;    Blue = 8'h3e;
end 12'hc5d:    begin Red = 8'h0c;    Green = 8'h87;    Blue = 8'hae;
end 12'hc5e:    begin Red = 8'h0c;    Green = 8'h76;    Blue = 8'he3;
end 12'hc5f:    begin Red = 8'hdb;    Green = 8'h99;    Blue = 8'hc8;
end 12'hc60:    begin Red = 8'h87;    Green = 8'h5e;    Blue = 8'h7e;
end 12'hc61:    begin Red = 8'h9e;    Green = 8'h6d;    Blue = 8'h93;
end 12'hc62:    begin Red = 8'h80;    Green = 8'h56;    Blue = 8'h71;
end 12'hc63:    begin Red = 8'h9b;    Green = 8'h88;    Blue = 8'h3a;
end 12'hc64:    begin Red = 8'hb7;    Green = 8'h8d;    Blue = 8'h45;
end 12'hc65:    begin Red = 8'ha8;    Green = 8'h8c;    Blue = 8'h35;
end 12'hc66:    begin Red = 8'hb1;    Green = 8'h8d;    Blue = 8'h45;
end 12'hc67:    begin Red = 8'hbc;    Green = 8'h86;    Blue = 8'h41;
end 12'hc68:    begin Red = 8'hfc;    Green = 8'he9;    Blue = 8'haa;
end 12'hc69:    begin Red = 8'hc7;    Green = 8'h90;    Blue = 8'hba;
end 12'hc6a:    begin Red = 8'hff;    Green = 8'hfc;    Blue = 8'hd7;
end 12'hc6b:    begin Red = 8'hb1;    Green = 8'h87;    Blue = 8'h26;
end 12'hc6c:    begin Red = 8'h79;    Green = 8'h6a;    Blue = 8'h2c;
end 12'hc6d:    begin Red = 8'hae;    Green = 8'h95;    Blue = 8'h62;
end 12'hc6e:    begin Red = 8'h0c;    Green = 8'h77;    Blue = 8'had;
end 12'hc6f:    begin Red = 8'h64;    Green = 8'h3e;    Blue = 8'h5d;
end 12'hc70:    begin Red = 8'h81;    Green = 8'h49;    Blue = 8'h6e;
end 12'hc71:    begin Red = 8'h62;    Green = 8'h3a;    Blue = 8'h57;
end 12'hc72:    begin Red = 8'h94;    Green = 8'h68;    Blue = 8'h92;
end 12'hc73:    begin Red = 8'h58;    Green = 8'h56;    Blue = 8'h50;
end 12'hc74:    begin Red = 8'h48;    Green = 8'h52;    Blue = 8'h4c;
end 12'hc75:    begin Red = 8'h4d;    Green = 8'h51;    Blue = 8'h49;
end 12'hc76:    begin Red = 8'hff;    Green = 8'hf4;    Blue = 8'hb3;
end 12'hc77:    begin Red = 8'h7c;    Green = 8'h47;    Blue = 8'h6b;
end 12'hc78:    begin Red = 8'hb9;    Green = 8'h97;    Blue = 8'h40;
end 12'hc79:    begin Red = 8'hc3;    Green = 8'h99;    Blue = 8'h50;
end 12'hc7a:    begin Red = 8'h9c;    Green = 8'ha7;    Blue = 8'h3e;
end 12'hc7b:    begin Red = 8'h7f;    Green = 8'h69;    Blue = 8'h2a;
end 12'hc7c:    begin Red = 8'h52;    Green = 8'h4d;    Blue = 8'h2a;
end 12'hc7d:    begin Red = 8'h0f;    Green = 8'h38;    Blue = 8'hb0;
end 12'hc7e:    begin Red = 8'h0f;    Green = 8'h39;    Blue = 8'h3e;
end 12'hc7f:    begin Red = 8'h89;    Green = 8'h78;    Blue = 8'h3c;
end 12'hc80:    begin Red = 8'h84;    Green = 8'h77;    Blue = 8'h3a;
end 12'hc81:    begin Red = 8'ha5;    Green = 8'h8f;    Blue = 8'h4f;
end 12'hc82:    begin Red = 8'h5e;    Green = 8'h54;    Blue = 8'h55;
end 12'hc83:    begin Red = 8'h52;    Green = 8'h4f;    Blue = 8'h5a;
end 12'hc84:    begin Red = 8'h5a;    Green = 8'h56;    Blue = 8'h5f;
end 12'hc85:    begin Red = 8'h42;    Green = 8'h4f;    Blue = 8'h4e;
end 12'hc86:    begin Red = 8'hab;    Green = 8'h6a;    Blue = 8'ha1;
end 12'hc87:    begin Red = 8'hb4;    Green = 8'h6b;    Blue = 8'h99;
end 12'hc88:    begin Red = 8'h60;    Green = 8'h5f;    Blue = 8'h55;
end 12'hc89:    begin Red = 8'h89;    Green = 8'h4f;    Blue = 8'h7f;
end 12'hc8a:    begin Red = 8'h87;    Green = 8'h64;    Blue = 8'h1c;
end 12'hc8b:    begin Red = 8'h08;    Green = 8'h38;    Blue = 8'h90;
end 12'hc8c:    begin Red = 8'h7e;    Green = 8'h6e;    Blue = 8'h29;
end 12'hc8d:    begin Red = 8'h0f;    Green = 8'hb8;    Blue = 8'h90;
end 12'hc8e:    begin Red = 8'h0f;    Green = 8'h59;    Blue = 8'h10;
end 12'hc8f:    begin Red = 8'h0e;    Green = 8'h69;    Blue = 8'h1e;
end 12'hc90:    begin Red = 8'h0f;    Green = 8'h09;    Blue = 8'h7e;
end 12'hc91:    begin Red = 8'h0c;    Green = 8'h87;    Blue = 8'h9b;
end 12'hc92:    begin Red = 8'hc2;    Green = 8'h77;    Blue = 8'h14;
end 12'hc93:    begin Red = 8'h0b;    Green = 8'he6;    Blue = 8'hf1;
end 12'hc94:    begin Red = 8'ha9;    Green = 8'h91;    Blue = 8'h57;
end 12'hc95:    begin Red = 8'hff;    Green = 8'hd9;    Blue = 8'h92;
end 12'hc96:    begin Red = 8'hfe;    Green = 8'hcf;    Blue = 8'h88;
end 12'hc97:    begin Red = 8'hd6;    Green = 8'h9f;    Blue = 8'h58;
end 12'hc98:    begin Red = 8'hc9;    Green = 8'ha3;    Blue = 8'h64;
end 12'hc99:    begin Red = 8'he4;    Green = 8'hb6;    Blue = 8'h6d;
end 12'hc9a:    begin Red = 8'ha0;    Green = 8'hab;    Blue = 8'h71;
end 12'hc9b:    begin Red = 8'h85;    Green = 8'h71;    Blue = 8'h35;
end 12'hc9c:    begin Red = 8'h42;    Green = 8'h58;    Blue = 8'h50;
end 12'hc9d:    begin Red = 8'h90;    Green = 8'h94;    Blue = 8'h66;
end 12'hc9e:    begin Red = 8'h9e;    Green = 8'h66;    Blue = 8'h89;
end 12'hc9f:    begin Red = 8'h96;    Green = 8'h9c;    Blue = 8'h2d;
end 12'hca0:    begin Red = 8'h78;    Green = 8'h6c;    Blue = 8'h33;
end 12'hca1:    begin Red = 8'ha8;    Green = 8'hb9;    Blue = 8'h80;
end 12'hca2:    begin Red = 8'hf6;    Green = 8'h9a;    Blue = 8'h11;
end 12'hca3:    begin Red = 8'hf4;    Green = 8'h97;    Blue = 8'h16;
end 12'hca4:    begin Red = 8'hf8;    Green = 8'h92;    Blue = 8'h17;
end 12'hca5:    begin Red = 8'h0b;    Green = 8'hd7;    Blue = 8'h7f;
end 12'hca6:    begin Red = 8'h0c;    Green = 8'h77;    Blue = 8'h8d;
end 12'hca7:    begin Red = 8'h0c;    Green = 8'h37;    Blue = 8'h01;
end 12'hca8:    begin Red = 8'hcc;    Green = 8'ha7;    Blue = 8'h6f;
end 12'hca9:    begin Red = 8'hbf;    Green = 8'h99;    Blue = 8'h67;
end 12'hcaa:    begin Red = 8'h96;    Green = 8'h9a;    Blue = 8'h36;
end 12'hcab:    begin Red = 8'h0f;    Green = 8'h19;    Blue = 8'h49;
end 12'hcac:    begin Red = 8'h0f;    Green = 8'hea;    Blue = 8'h5a;
end 12'hcad:    begin Red = 8'h0f;    Green = 8'hea;    Blue = 8'h33;
end 12'hcae:    begin Red = 8'hf1;    Green = 8'h91;    Blue = 8'h16;
end 12'hcaf:    begin Red = 8'h0d;    Green = 8'ha8;    Blue = 8'h48;
end 12'hcb0:    begin Red = 8'hc6;    Green = 8'h7e;    Blue = 8'h12;
end 12'hcb1:    begin Red = 8'he2;    Green = 8'hae;    Blue = 8'h6f;
end 12'hcb2:    begin Red = 8'h01;    Green = 8'h3d;    Blue = 8'h18;
end 12'hcb3:    begin Red = 8'h11;    Green = 8'h10;    Blue = 8'h17;
end 12'hcb4:    begin Red = 8'h24;    Green = 8'h1e;    Blue = 8'h2b;
end 12'hcb5:    begin Red = 8'hea;    Green = 8'he6;    Blue = 8'hc3;
end 12'hcb6:    begin Red = 8'h7a;    Green = 8'h3d;    Blue = 8'h1b;
end 12'hcb7:    begin Red = 8'h78;    Green = 8'h62;    Blue = 8'h2c;
end 12'hcb8:    begin Red = 8'h53;    Green = 8'h46;    Blue = 8'h35;
end 12'hcb9:    begin Red = 8'h2f;    Green = 8'h2a;    Blue = 8'h26;
end 12'hcba:    begin Red = 8'h00;    Green = 8'hfc;    Blue = 8'h16;
end 12'hcbb:    begin Red = 8'he6;    Green = 8'he2;    Blue = 8'hca;
end 12'hcbc:    begin Red = 8'ha7;    Green = 8'ha4;    Blue = 8'h74;
end 12'hcbd:    begin Red = 8'haa;    Green = 8'h7f;    Blue = 8'h4d;
end 12'hcbe:    begin Red = 8'h00;    Green = 8'h05;    Blue = 8'h05;
end 12'hcbf:    begin Red = 8'h01;    Green = 8'h5f;    Blue = 8'h12;
end 12'hcc0:    begin Red = 8'h34;    Green = 8'h22;    Blue = 8'h17;
end 12'hcc1:    begin Red = 8'h35;    Green = 8'h1d;    Blue = 8'h18;
end 12'hcc2:    begin Red = 8'h00;    Green = 8'h01;    Blue = 8'h32;
end 12'hcc3:    begin Red = 8'h53;    Green = 8'h4e;    Blue = 8'h4d;
end 12'hcc4:    begin Red = 8'h1a;    Green = 8'h10;    Blue = 8'h18;
end 12'hcc5:    begin Red = 8'he1;    Green = 8'hc9;    Blue = 8'hae;
end 12'hcc6:    begin Red = 8'h9d;    Green = 8'h97;    Blue = 8'h4d;
end 12'hcc7:    begin Red = 8'h4b;    Green = 8'h4b;    Blue = 8'h4b;
end 12'hcc8:    begin Red = 8'he3;    Green = 8'hd8;    Blue = 8'hb3;
end 12'hcc9:    begin Red = 8'had;    Green = 8'hb0;    Blue = 8'h78;
end 12'hcca:    begin Red = 8'h5a;    Green = 8'h41;    Blue = 8'h15;
end 12'hccb:    begin Red = 8'h05;    Green = 8'he3;    Blue = 8'h84;
end 12'hccc:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'h29;
end 12'hccd:    begin Red = 8'h07;    Green = 8'he4;    Blue = 8'heb;
end 12'hcce:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'hfc;
end 12'hccf:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h25;
end 12'hcd0:    begin Red = 8'h05;    Green = 8'h83;    Blue = 8'h29;
end 12'hcd1:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'h6d;
end 12'hcd2:    begin Red = 8'h07;    Green = 8'h34;    Blue = 8'h5e;
end 12'hcd3:    begin Red = 8'h07;    Green = 8'h14;    Blue = 8'h3b;
end 12'hcd4:    begin Red = 8'he1;    Green = 8'hed;    Blue = 8'hc2;
end 12'hcd5:    begin Red = 8'h67;    Green = 8'h46;    Blue = 8'h15;
end 12'hcd6:    begin Red = 8'h88;    Green = 8'h8d;    Blue = 8'h6c;
end 12'hcd7:    begin Red = 8'ha0;    Green = 8'h8e;    Blue = 8'h75;
end 12'hcd8:    begin Red = 8'h00;    Green = 8'h0a;    Blue = 8'h46;
end 12'hcd9:    begin Red = 8'h02;    Green = 8'h91;    Blue = 8'hec;
end 12'hcda:    begin Red = 8'h30;    Green = 8'h1b;    Blue = 8'h15;
end 12'hcdb:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'hbb;
end 12'hcdc:    begin Red = 8'h02;    Green = 8'h31;    Blue = 8'he1;
end 12'hcdd:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'hdd;
end 12'hcde:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'hfe;
end 12'hcdf:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'hca;
end 12'hce0:    begin Red = 8'h47;    Green = 8'h4d;    Blue = 8'h53;
end 12'hce1:    begin Red = 8'h2b;    Green = 8'h34;    Blue = 8'h4d;
end 12'hce2:    begin Red = 8'h33;    Green = 8'h39;    Blue = 8'h53;
end 12'hce3:    begin Red = 8'h5b;    Green = 8'h5b;    Blue = 8'h4b;
end 12'hce4:    begin Red = 8'h82;    Green = 8'h81;    Blue = 8'h4b;
end 12'hce5:    begin Red = 8'hcc;    Green = 8'hd6;    Blue = 8'hba;
end 12'hce6:    begin Red = 8'hf9;    Green = 8'hec;    Blue = 8'hdd;
end 12'hce7:    begin Red = 8'h2c;    Green = 8'h21;    Blue = 8'h24;
end 12'hce8:    begin Red = 8'h01;    Green = 8'h6b;    Blue = 8'h10;
end 12'hce9:    begin Red = 8'h9e;    Green = 8'h9c;    Blue = 8'h38;
end 12'hcea:    begin Red = 8'h33;    Green = 8'h31;    Blue = 8'h4e;
end 12'hceb:    begin Red = 8'h3c;    Green = 8'h38;    Blue = 8'h51;
end 12'hcec:    begin Red = 8'h56;    Green = 8'h5d;    Blue = 8'h4c;
end 12'hced:    begin Red = 8'hd6;    Green = 8'hc1;    Blue = 8'h9e;
end 12'hcee:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'hb2;
end 12'hcef:    begin Red = 8'h04;    Green = 8'h62;    Blue = 8'h50;
end 12'hcf0:    begin Red = 8'h02;    Green = 8'h81;    Blue = 8'h80;
end 12'hcf1:    begin Red = 8'h04;    Green = 8'h01;    Blue = 8'he3;
end 12'hcf2:    begin Red = 8'h08;    Green = 8'h75;    Blue = 8'h1c;
end 12'hcf3:    begin Red = 8'h08;    Green = 8'h45;    Blue = 8'h0f;
end 12'hcf4:    begin Red = 8'h08;    Green = 8'h55;    Blue = 8'h1f;
end 12'hcf5:    begin Red = 8'h08;    Green = 8'h35;    Blue = 8'h2b;
end 12'hcf6:    begin Red = 8'h05;    Green = 8'h63;    Blue = 8'h5d;
end 12'hcf7:    begin Red = 8'h05;    Green = 8'h63;    Blue = 8'h36;
end 12'hcf8:    begin Red = 8'h07;    Green = 8'hd4;    Blue = 8'hcd;
end 12'hcf9:    begin Red = 8'h07;    Green = 8'h04;    Blue = 8'h7b;
end 12'hcfa:    begin Red = 8'hd8;    Green = 8'he5;    Blue = 8'hbd;
end 12'hcfb:    begin Red = 8'h06;    Green = 8'ha4;    Blue = 8'h15;
end 12'hcfc:    begin Red = 8'h06;    Green = 8'h23;    Blue = 8'hc8;
end 12'hcfd:    begin Red = 8'h8b;    Green = 8'h67;    Blue = 8'h16;
end 12'hcfe:    begin Red = 8'h92;    Green = 8'h66;    Blue = 8'h18;
end 12'hcff:    begin Red = 8'h85;    Green = 8'h6a;    Blue = 8'h16;
end 12'hd00:    begin Red = 8'h8a;    Green = 8'h6a;    Blue = 8'h10;
end 12'hd01:    begin Red = 8'h07;    Green = 8'hf6;    Blue = 8'hb5;
end 12'hd02:    begin Red = 8'h08;    Green = 8'h46;    Blue = 8'h26;
end 12'hd03:    begin Red = 8'h4c;    Green = 8'h33;    Blue = 8'h32;
end 12'hd04:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h6f;
end 12'hd05:    begin Red = 8'h48;    Green = 8'h2d;    Blue = 8'h32;
end 12'hd06:    begin Red = 8'h71;    Green = 8'h3c;    Blue = 8'h61;
end 12'hd07:    begin Red = 8'h5d;    Green = 8'h36;    Blue = 8'h59;
end 12'hd08:    begin Red = 8'h00;    Green = 8'h13;    Blue = 8'h0d;
end 12'hd09:    begin Red = 8'h2d;    Green = 8'h2d;    Blue = 8'h31;
end 12'hd0a:    begin Red = 8'h52;    Green = 8'h4d;    Blue = 8'h48;
end 12'hd0b:    begin Red = 8'h00;    Green = 8'h95;    Blue = 8'h1b;
end 12'hd0c:    begin Red = 8'hd3;    Green = 8'ha5;    Blue = 8'h23;
end 12'hd0d:    begin Red = 8'hb9;    Green = 8'h3f;    Blue = 8'h36;
end 12'hd0e:    begin Red = 8'hc5;    Green = 8'ha5;    Blue = 8'h4e;
end 12'hd0f:    begin Red = 8'hbf;    Green = 8'h95;    Blue = 8'h40;
end 12'hd10:    begin Red = 8'h01;    Green = 8'h3c;    Blue = 8'h12;
end 12'hd11:    begin Red = 8'h2f;    Green = 8'h25;    Blue = 8'h2c;
end 12'hd12:    begin Red = 8'h01;    Green = 8'h6c;    Blue = 8'h16;
end 12'hd13:    begin Red = 8'h99;    Green = 8'h9d;    Blue = 8'h3d;
end 12'hd14:    begin Red = 8'h81;    Green = 8'h6e;    Blue = 8'h2f;
end 12'hd15:    begin Red = 8'h02;    Green = 8'hf1;    Blue = 8'h40;
end 12'hd16:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'hd1;
end 12'hd17:    begin Red = 8'h06;    Green = 8'hb4;    Blue = 8'h28;
end 12'hd18:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'he4;
end 12'hd19:    begin Red = 8'h06;    Green = 8'hd4;    Blue = 8'h04;
end 12'hd1a:    begin Red = 8'h06;    Green = 8'hc3;    Blue = 8'hf3;
end 12'hd1b:    begin Red = 8'h06;    Green = 8'ha3;    Blue = 8'hf6;
end 12'hd1c:    begin Red = 8'h06;    Green = 8'h84;    Blue = 8'h06;
end 12'hd1d:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'he4;
end 12'hd1e:    begin Red = 8'h04;    Green = 8'h42;    Blue = 8'h81;
end 12'hd1f:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h60;
end 12'hd20:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h91;
end 12'hd21:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'he9;
end 12'hd22:    begin Red = 8'h05;    Green = 8'hd3;    Blue = 8'hc4;
end 12'hd23:    begin Red = 8'h05;    Green = 8'h93;    Blue = 8'h73;
end 12'hd24:    begin Red = 8'h05;    Green = 8'h73;    Blue = 8'h48;
end 12'hd25:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h15;
end 12'hd26:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h46;
end 12'hd27:    begin Red = 8'h05;    Green = 8'h33;    Blue = 8'h04;
end 12'hd28:    begin Red = 8'h33;    Green = 8'h3f;    Blue = 8'h71;
end 12'hd29:    begin Red = 8'h30;    Green = 8'h45;    Blue = 8'h6b;
end 12'hd2a:    begin Red = 8'h50;    Green = 8'h39;    Blue = 8'h3a;
end 12'hd2b:    begin Red = 8'h4e;    Green = 8'h31;    Blue = 8'h3e;
end 12'hd2c:    begin Red = 8'h55;    Green = 8'h3b;    Blue = 8'h40;
end 12'hd2d:    begin Red = 8'h4b;    Green = 8'h37;    Blue = 8'h3a;
end 12'hd2e:    begin Red = 8'h53;    Green = 8'h37;    Blue = 8'h47;
end 12'hd2f:    begin Red = 8'h02;    Green = 8'h2b;    Blue = 8'h24;
end 12'hd30:    begin Red = 8'hf0;    Green = 8'he8;    Blue = 8'hce;
end 12'hd31:    begin Red = 8'hbc;    Green = 8'ha7;    Blue = 8'h4a;
end 12'hd32:    begin Red = 8'hf2;    Green = 8'he8;    Blue = 8'hdd;
end 12'hd33:    begin Red = 8'h00;    Green = 8'h2d;    Blue = 8'h62;
end 12'hd34:    begin Red = 8'h0e;    Green = 8'h38;    Blue = 8'h59;
end 12'hd35:    begin Red = 8'h51;    Green = 8'hc0;    Blue = 8'hf6;
end 12'hd36:    begin Red = 8'hd7;    Green = 8'hfc;    Blue = 8'hf6;
end 12'hd37:    begin Red = 8'hd6;    Green = 8'hfb;    Blue = 8'hed;
end 12'hd38:    begin Red = 8'hbf;    Green = 8'h53;    Blue = 8'h57;
end 12'hd39:    begin Red = 8'ha1;    Green = 8'ha2;    Blue = 8'h6b;
end 12'hd3a:    begin Red = 8'h88;    Green = 8'h8f;    Blue = 8'h5f;
end 12'hd3b:    begin Red = 8'h72;    Green = 8'h7c;    Blue = 8'h41;
end 12'hd3c:    begin Red = 8'h06;    Green = 8'h83;    Blue = 8'h51;
end 12'hd3d:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'h77;
end 12'hd3e:    begin Red = 8'h99;    Green = 8'h98;    Blue = 8'h6a;
end 12'hd3f:    begin Red = 8'h8e;    Green = 8'h8d;    Blue = 8'h60;
end 12'hd40:    begin Red = 8'hb4;    Green = 8'hbd;    Blue = 8'h92;
end 12'hd41:    begin Red = 8'h4d;    Green = 8'h5e;    Blue = 8'h35;
end 12'hd42:    begin Red = 8'h15;    Green = 8'h2b;    Blue = 8'h37;
end 12'hd43:    begin Red = 8'h17;    Green = 8'h29;    Blue = 8'h3d;
end 12'hd44:    begin Red = 8'h2d;    Green = 8'h2d;    Blue = 8'h45;
end 12'hd45:    begin Red = 8'h3f;    Green = 8'h4e;    Blue = 8'h5b;
end 12'hd46:    begin Red = 8'h3f;    Green = 8'h44;    Blue = 8'h50;
end 12'hd47:    begin Red = 8'h3d;    Green = 8'h3f;    Blue = 8'h4e;
end 12'hd48:    begin Red = 8'h3a;    Green = 8'h48;    Blue = 8'h5d;
end 12'hd49:    begin Red = 8'h08;    Green = 8'h26;    Blue = 8'h26;
end 12'hd4a:    begin Red = 8'had;    Green = 8'h92;    Blue = 8'h7c;
end 12'hd4b:    begin Red = 8'hd0;    Green = 8'hb5;    Blue = 8'h7b;
end 12'hd4c:    begin Red = 8'hfe;    Green = 8'hf9;    Blue = 8'hbc;
end 12'hd4d:    begin Red = 8'h4f;    Green = 8'h37;    Blue = 8'h40;
end 12'hd4e:    begin Red = 8'h5d;    Green = 8'h3a;    Blue = 8'h47;
end 12'hd4f:    begin Red = 8'h4d;    Green = 8'h3d;    Blue = 8'h41;
end 12'hd50:    begin Red = 8'h47;    Green = 8'h2c;    Blue = 8'h39;
end 12'hd51:    begin Red = 8'h52;    Green = 8'h32;    Blue = 8'h43;
end 12'hd52:    begin Red = 8'h43;    Green = 8'h2c;    Blue = 8'h3e;
end 12'hd53:    begin Red = 8'h02;    Green = 8'h01;    Blue = 8'h76;
end 12'hd54:    begin Red = 8'hb6;    Green = 8'h3f;    Blue = 8'h3c;
end 12'hd55:    begin Red = 8'hb6;    Green = 8'h3f;    Blue = 8'h30;
end 12'hd56:    begin Red = 8'hbd;    Green = 8'hae;    Blue = 8'h48;
end 12'hd57:    begin Red = 8'hac;    Green = 8'h81;    Blue = 8'h2b;
end 12'hd58:    begin Red = 8'h2b;    Green = 8'h5b;    Blue = 8'h76;
end 12'hd59:    begin Red = 8'h33;    Green = 8'h5a;    Blue = 8'h7a;
end 12'hd5a:    begin Red = 8'h1e;    Green = 8'h5f;    Blue = 8'h74;
end 12'hd5b:    begin Red = 8'h50;    Green = 8'hce;    Blue = 8'heb;
end 12'hd5c:    begin Red = 8'h52;    Green = 8'ha1;    Blue = 8'hd3;
end 12'hd5d:    begin Red = 8'h4f;    Green = 8'hab;    Blue = 8'he5;
end 12'hd5e:    begin Red = 8'hd5;    Green = 8'h4f;    Blue = 8'h3d;
end 12'hd5f:    begin Red = 8'he9;    Green = 8'heb;    Blue = 8'hb2;
end 12'hd60:    begin Red = 8'h83;    Green = 8'h74;    Blue = 8'h29;
end 12'hd61:    begin Red = 8'h00;    Green = 8'h00;    Blue = 8'h18;
end 12'hd62:    begin Red = 8'h00;    Green = 8'h78;    Blue = 8'h19;
end 12'hd63:    begin Red = 8'h2c;    Green = 8'h30;    Blue = 8'h2a;
end 12'hd64:    begin Red = 8'hba;    Green = 8'ha8;    Blue = 8'h95;
end 12'hd65:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'hd2;
end 12'hd66:    begin Red = 8'h9c;    Green = 8'h92;    Blue = 8'h62;
end 12'hd67:    begin Red = 8'h97;    Green = 8'h90;    Blue = 8'h58;
end 12'hd68:    begin Red = 8'h98;    Green = 8'h90;    Blue = 8'h5d;
end 12'hd69:    begin Red = 8'h8b;    Green = 8'h87;    Blue = 8'h52;
end 12'hd6a:    begin Red = 8'h90;    Green = 8'h87;    Blue = 8'h52;
end 12'hd6b:    begin Red = 8'h85;    Green = 8'h82;    Blue = 8'h50;
end 12'hd6c:    begin Red = 8'h7f;    Green = 8'h7d;    Blue = 8'h43;
end 12'hd6d:    begin Red = 8'h71;    Green = 8'h75;    Blue = 8'h3c;
end 12'hd6e:    begin Red = 8'h06;    Green = 8'h13;    Blue = 8'hc3;
end 12'hd6f:    begin Red = 8'ha4;    Green = 8'haf;    Blue = 8'h81;
end 12'hd70:    begin Red = 8'h52;    Green = 8'h56;    Blue = 8'h2c;
end 12'hd71:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h78;
end 12'hd72:    begin Red = 8'hac;    Green = 8'h88;    Blue = 8'h57;
end 12'hd73:    begin Red = 8'h81;    Green = 8'hcf;    Blue = 8'hc7;
end 12'hd74:    begin Red = 8'h4c;    Green = 8'h8d;    Blue = 8'ha3;
end 12'hd75:    begin Red = 8'h48;    Green = 8'h7d;    Blue = 8'h93;
end 12'hd76:    begin Red = 8'h46;    Green = 8'h44;    Blue = 8'h50;
end 12'hd77:    begin Red = 8'h37;    Green = 8'h41;    Blue = 8'h44;
end 12'hd78:    begin Red = 8'h51;    Green = 8'h7e;    Blue = 8'h94;
end 12'hd79:    begin Red = 8'h2f;    Green = 8'h18;    Blue = 8'h29;
end 12'hd7a:    begin Red = 8'h29;    Green = 8'h18;    Blue = 8'h27;
end 12'hd7b:    begin Red = 8'h40;    Green = 8'h26;    Blue = 8'h2f;
end 12'hd7c:    begin Red = 8'h38;    Green = 8'h21;    Blue = 8'h26;
end 12'hd7d:    begin Red = 8'h3a;    Green = 8'h28;    Blue = 8'h23;
end 12'hd7e:    begin Red = 8'h01;    Green = 8'hf1;    Blue = 8'h59;
end 12'hd7f:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'h11;
end 12'hd80:    begin Red = 8'h4a;    Green = 8'h28;    Blue = 8'h28;
end 12'hd81:    begin Red = 8'h79;    Green = 8'h47;    Blue = 8'h42;
end 12'hd82:    begin Red = 8'h2d;    Green = 8'h19;    Blue = 8'h1a;
end 12'hd83:    begin Red = 8'h5d;    Green = 8'h4b;    Blue = 8'h59;
end 12'hd84:    begin Red = 8'h45;    Green = 8'h2c;    Blue = 8'h2d;
end 12'hd85:    begin Red = 8'h63;    Green = 8'h4e;    Blue = 8'h57;
end 12'hd86:    begin Red = 8'h00;    Green = 8'h0b;    Blue = 8'h19;
end 12'hd87:    begin Red = 8'h2d;    Green = 8'h3b;    Blue = 8'h50;
end 12'hd88:    begin Red = 8'h1e;    Green = 8'h4d;    Blue = 8'h61;
end 12'hd89:    begin Red = 8'h02;    Green = 8'h31;    Blue = 8'h17;
end 12'hd8a:    begin Red = 8'h34;    Green = 8'h2d;    Blue = 8'h32;
end 12'hd8b:    begin Red = 8'h52;    Green = 8'ha1;    Blue = 8'hdc;
end 12'hd8c:    begin Red = 8'h4e;    Green = 8'ha7;    Blue = 8'hd8;
end 12'hd8d:    begin Red = 8'h99;    Green = 8'h98;    Blue = 8'h3b;
end 12'hd8e:    begin Red = 8'h77;    Green = 8'h69;    Blue = 8'h25;
end 12'hd8f:    begin Red = 8'ha0;    Green = 8'ha7;    Blue = 8'h7a;
end 12'hd90:    begin Red = 8'he3;    Green = 8'hbe;    Blue = 8'h83;
end 12'hd91:    begin Red = 8'h00;    Green = 8'h2c;    Blue = 8'he3;
end 12'hd92:    begin Red = 8'h9f;    Green = 8'h98;    Blue = 8'h60;
end 12'hd93:    begin Red = 8'h68;    Green = 8'h6e;    Blue = 8'h3a;
end 12'hd94:    begin Red = 8'h6e;    Green = 8'h6f;    Blue = 8'h3d;
end 12'hd95:    begin Red = 8'h85;    Green = 8'h7b;    Blue = 8'h4e;
end 12'hd96:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h89;
end 12'hd97:    begin Red = 8'h5b;    Green = 8'hc3;    Blue = 8'hba;
end 12'hd98:    begin Red = 8'h69;    Green = 8'hc7;    Blue = 8'hc0;
end 12'hd99:    begin Red = 8'h4e;    Green = 8'h88;    Blue = 8'ha9;
end 12'hd9a:    begin Red = 8'h53;    Green = 8'h8f;    Blue = 8'ha0;
end 12'hd9b:    begin Red = 8'h5a;    Green = 8'h8c;    Blue = 8'haf;
end 12'hd9c:    begin Red = 8'h48;    Green = 8'h78;    Blue = 8'h92;
end 12'hd9d:    begin Red = 8'h39;    Green = 8'h74;    Blue = 8'h8c;
end 12'hd9e:    begin Red = 8'hc5;    Green = 8'hb0;    Blue = 8'h74;
end 12'hd9f:    begin Red = 8'h2c;    Green = 8'h16;    Blue = 8'h22;
end 12'hda0:    begin Red = 8'h7b;    Green = 8'h46;    Blue = 8'h48;
end 12'hda1:    begin Red = 8'h5e;    Green = 8'h51;    Blue = 8'h5b;
end 12'hda2:    begin Red = 8'h5c;    Green = 8'h4e;    Blue = 8'h53;
end 12'hda3:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h38;
end 12'hda4:    begin Red = 8'h63;    Green = 8'h53;    Blue = 8'h58;
end 12'hda5:    begin Red = 8'h67;    Green = 8'h59;    Blue = 8'h61;
end 12'hda6:    begin Red = 8'hfc;    Green = 8'hc1;    Blue = 8'h2a;
end 12'hda7:    begin Red = 8'h42;    Green = 8'h42;    Blue = 8'h55;
end 12'hda8:    begin Red = 8'hc6;    Green = 8'h3b;    Blue = 8'h30;
end 12'hda9:    begin Red = 8'had;    Green = 8'h1d;    Blue = 8'h13;
end 12'hdaa:    begin Red = 8'ha8;    Green = 8'h8e;    Blue = 8'h2e;
end 12'hdab:    begin Red = 8'h34;    Green = 8'h4c;    Blue = 8'h71;
end 12'hdac:    begin Red = 8'h51;    Green = 8'hb2;    Blue = 8'hed;
end 12'hdad:    begin Red = 8'h54;    Green = 8'hc6;    Blue = 8'hf6;
end 12'hdae:    begin Red = 8'h4d;    Green = 8'hb2;    Blue = 8'he7;
end 12'hdaf:    begin Red = 8'h03;    Green = 8'h21;    Blue = 8'h57;
end 12'hdb0:    begin Red = 8'h52;    Green = 8'ha8;    Blue = 8'hec;
end 12'hdb1:    begin Red = 8'haa;    Green = 8'hac;    Blue = 8'h3b;
end 12'hdb2:    begin Red = 8'hf2;    Green = 8'hbb;    Blue = 8'h22;
end 12'hdb3:    begin Red = 8'hf9;    Green = 8'hbf;    Blue = 8'h25;
end 12'hdb4:    begin Red = 8'h53;    Green = 8'h53;    Blue = 8'h4c;
end 12'hdb5:    begin Red = 8'h36;    Green = 8'h36;    Blue = 8'h3a;
end 12'hdb6:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h21;
end 12'hdb7:    begin Red = 8'h04;    Green = 8'ha2;    Blue = 8'hd0;
end 12'hdb8:    begin Red = 8'h7a;    Green = 8'h79;    Blue = 8'h46;
end 12'hdb9:    begin Red = 8'h80;    Green = 8'h79;    Blue = 8'h48;
end 12'hdba:    begin Red = 8'h85;    Green = 8'hce;    Blue = 8'hcf;
end 12'hdbb:    begin Red = 8'h95;    Green = 8'he8;    Blue = 8'he2;
end 12'hdbc:    begin Red = 8'h95;    Green = 8'he7;    Blue = 8'he7;
end 12'hdbd:    begin Red = 8'h32;    Green = 8'h1e;    Blue = 8'h29;
end 12'hdbe:    begin Red = 8'h3e;    Green = 8'h26;    Blue = 8'h34;
end 12'hdbf:    begin Red = 8'h77;    Green = 8'h41;    Blue = 8'h48;
end 12'hdc0:    begin Red = 8'h3a;    Green = 8'h23;    Blue = 8'h2b;
end 12'hdc1:    begin Red = 8'h50;    Green = 8'h42;    Blue = 8'h4a;
end 12'hdc2:    begin Red = 8'h27;    Green = 8'h25;    Blue = 8'h27;
end 12'hdc3:    begin Red = 8'hb9;    Green = 8'h94;    Blue = 8'h4f;
end 12'hdc4:    begin Red = 8'h40;    Green = 8'h68;    Blue = 8'h81;
end 12'hdc5:    begin Red = 8'h48;    Green = 8'h7d;    Blue = 8'h9d;
end 12'hdc6:    begin Red = 8'h25;    Green = 8'h16;    Blue = 8'h1c;
end 12'hdc7:    begin Red = 8'h00;    Green = 8'h1e;    Blue = 8'h30;
end 12'hdc8:    begin Red = 8'h40;    Green = 8'h67;    Blue = 8'h87;
end 12'hdc9:    begin Red = 8'h51;    Green = 8'had;    Blue = 8'hed;
end 12'hdca:    begin Red = 8'h47;    Green = 8'ha2;    Blue = 8'hd9;
end 12'hdcb:    begin Red = 8'hcd;    Green = 8'ha6;    Blue = 8'h25;
end 12'hdcc:    begin Red = 8'h00;    Green = 8'hb9;    Blue = 8'h20;
end 12'hdcd:    begin Red = 8'h75;    Green = 8'h71;    Blue = 8'h43;
end 12'hdce:    begin Red = 8'h57;    Green = 8'h55;    Blue = 8'h58;
end 12'hdcf:    begin Red = 8'hb8;    Green = 8'hd9;    Blue = 8'hce;
end 12'hdd0:    begin Red = 8'h7a;    Green = 8'hc5;    Blue = 8'hd0;
end 12'hdd1:    begin Red = 8'h8c;    Green = 8'hc9;    Blue = 8'hc9;
end 12'hdd2:    begin Red = 8'h82;    Green = 8'hca;    Blue = 8'hc8;
end 12'hdd3:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'h2e;
end 12'hdd4:    begin Red = 8'h35;    Green = 8'h25;    Blue = 8'h30;
end 12'hdd5:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'h3a;
end 12'hdd6:    begin Red = 8'h56;    Green = 8'hb7;    Blue = 8'hf4;
end 12'hdd7:    begin Red = 8'h2a;    Green = 8'h51;    Blue = 8'h67;
end 12'hdd8:    begin Red = 8'h41;    Green = 8'h6e;    Blue = 8'h84;
end 12'hdd9:    begin Red = 8'h3b;    Green = 8'h67;    Blue = 8'h84;
end 12'hdda:    begin Red = 8'h38;    Green = 8'h6f;    Blue = 8'h7b;
end 12'hddb:    begin Red = 8'h42;    Green = 8'h62;    Blue = 8'h87;
end 12'hddc:    begin Red = 8'h38;    Green = 8'h65;    Blue = 8'h7c;
end 12'hddd:    begin Red = 8'h3a;    Green = 8'h6e;    Blue = 8'h8c;
end 12'hdde:    begin Red = 8'hfb;    Green = 8'h4a;    Blue = 8'h21;
end 12'hddf:    begin Red = 8'hf1;    Green = 8'h54;    Blue = 8'h3a;
end 12'hde0:    begin Red = 8'h95;    Green = 8'h8b;    Blue = 8'h59;
end 12'hde1:    begin Red = 8'h8a;    Green = 8'h82;    Blue = 8'h54;
end 12'hde2:    begin Red = 8'h06;    Green = 8'h53;    Blue = 8'hf9;
end 12'hde3:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'hc3;
end 12'hde4:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h47;
end 12'hde5:    begin Red = 8'h48;    Green = 8'h3f;    Blue = 8'h48;
end 12'hde6:    begin Red = 8'h6e;    Green = 8'hcb;    Blue = 8'hc0;
end 12'hde7:    begin Red = 8'h79;    Green = 8'hc8;    Blue = 8'hc6;
end 12'hde8:    begin Red = 8'h74;    Green = 8'hcf;    Blue = 8'hd2;
end 12'hde9:    begin Red = 8'h73;    Green = 8'he3;    Blue = 8'he5;
end 12'hdea:    begin Red = 8'h74;    Green = 8'he6;    Blue = 8'heb;
end 12'hdeb:    begin Red = 8'h4d;    Green = 8'h2f;    Blue = 8'h44;
end 12'hdec:    begin Red = 8'hf3;    Green = 8'hfc;    Blue = 8'hc3;
end 12'hded:    begin Red = 8'h35;    Green = 8'h14;    Blue = 8'h24;
end 12'hdee:    begin Red = 8'h01;    Green = 8'h81;    Blue = 8'h30;
end 12'hdef:    begin Red = 8'h4c;    Green = 8'h31;    Blue = 8'h39;
end 12'hdf0:    begin Red = 8'h47;    Green = 8'h31;    Blue = 8'h37;
end 12'hdf1:    begin Red = 8'h01;    Green = 8'h36;    Blue = 8'h16;
end 12'hdf2:    begin Red = 8'h31;    Green = 8'h35;    Blue = 8'h3a;
end 12'hdf3:    begin Red = 8'h8d;    Green = 8'h7a;    Blue = 8'h69;
end 12'hdf4:    begin Red = 8'h5b;    Green = 8'hb8;    Blue = 8'hf2;
end 12'hdf5:    begin Red = 8'h5c;    Green = 8'hc4;    Blue = 8'hf6;
end 12'hdf6:    begin Red = 8'h29;    Green = 8'h4b;    Blue = 8'h5c;
end 12'hdf7:    begin Red = 8'h22;    Green = 8'h55;    Blue = 8'h60;
end 12'hdf8:    begin Red = 8'h33;    Green = 8'h5f;    Blue = 8'h7b;
end 12'hdf9:    begin Red = 8'h41;    Green = 8'h63;    Blue = 8'h80;
end 12'hdfa:    begin Red = 8'h35;    Green = 8'h6d;    Blue = 8'h84;
end 12'hdfb:    begin Red = 8'h3b;    Green = 8'h6e;    Blue = 8'h81;
end 12'hdfc:    begin Red = 8'h18;    Green = 8'h71;    Blue = 8'h92;
end 12'hdfd:    begin Red = 8'hff;    Green = 8'h38;    Blue = 8'h19;
end 12'hdfe:    begin Red = 8'hf9;    Green = 8'h30;    Blue = 8'h21;
end 12'hdff:    begin Red = 8'hae;    Green = 8'hb0;    Blue = 8'h42;
end 12'he00:    begin Red = 8'h58;    Green = 8'h4e;    Blue = 8'h25;
end 12'he01:    begin Red = 8'h3a;    Green = 8'h37;    Blue = 8'h41;
end 12'he02:    begin Red = 8'h9c;    Green = 8'ha2;    Blue = 8'h6f;
end 12'he03:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'hc4;
end 12'he04:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h35;
end 12'he05:    begin Red = 8'h84;    Green = 8'h91;    Blue = 8'h93;
end 12'he06:    begin Red = 8'h72;    Green = 8'h84;    Blue = 8'h87;
end 12'he07:    begin Red = 8'hb7;    Green = 8'hd8;    Blue = 8'hd7;
end 12'he08:    begin Red = 8'hb4;    Green = 8'hdc;    Blue = 8'hc9;
end 12'he09:    begin Red = 8'hbe;    Green = 8'hdf;    Blue = 8'hdd;
end 12'he0a:    begin Red = 8'hb2;    Green = 8'hef;    Blue = 8'hf3;
end 12'he0b:    begin Red = 8'hbd;    Green = 8'h63;    Blue = 8'h63;
end 12'he0c:    begin Red = 8'hbd;    Green = 8'h61;    Blue = 8'h5e;
end 12'he0d:    begin Red = 8'h08;    Green = 8'h46;    Blue = 8'h05;
end 12'he0e:    begin Red = 8'h3d;    Green = 8'h25;    Blue = 8'h39;
end 12'he0f:    begin Red = 8'h57;    Green = 8'h2c;    Blue = 8'h45;
end 12'he10:    begin Red = 8'he4;    Green = 8'hef;    Blue = 8'haf;
end 12'he11:    begin Red = 8'h48;    Green = 8'h2a;    Blue = 8'h40;
end 12'he12:    begin Red = 8'h3a;    Green = 8'h21;    Blue = 8'h32;
end 12'he13:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h02;
end 12'he14:    begin Red = 8'h00;    Green = 8'he2;    Blue = 8'h17;
end 12'he15:    begin Red = 8'h23;    Green = 8'h4f;    Blue = 8'h64;
end 12'he16:    begin Red = 8'h5c;    Green = 8'had;    Blue = 8'hf4;
end 12'he17:    begin Red = 8'h01;    Green = 8'h91;    Blue = 8'h00;
end 12'he18:    begin Red = 8'hea;    Green = 8'h4c;    Blue = 8'h3a;
end 12'he19:    begin Red = 8'hd8;    Green = 8'hf2;    Blue = 8'hcf;
end 12'he1a:    begin Red = 8'h04;    Green = 8'ha2;    Blue = 8'hd5;
end 12'he1b:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'h91;
end 12'he1c:    begin Red = 8'h45;    Green = 8'h48;    Blue = 8'h23;
end 12'he1d:    begin Red = 8'h8a;    Green = 8'h8c;    Blue = 8'h95;
end 12'he1e:    begin Red = 8'h7d;    Green = 8'h92;    Blue = 8'h95;
end 12'he1f:    begin Red = 8'h6b;    Green = 8'h81;    Blue = 8'h85;
end 12'he20:    begin Red = 8'hdc;    Green = 8'he4;    Blue = 8'hd9;
end 12'he21:    begin Red = 8'hb3;    Green = 8'hd6;    Blue = 8'hca;
end 12'he22:    begin Red = 8'hc1;    Green = 8'h36;    Blue = 8'h29;
end 12'he23:    begin Red = 8'hbd;    Green = 8'h4b;    Blue = 8'h46;
end 12'he24:    begin Red = 8'hbe;    Green = 8'h60;    Blue = 8'h57;
end 12'he25:    begin Red = 8'hb6;    Green = 8'h63;    Blue = 8'h56;
end 12'he26:    begin Red = 8'h4c;    Green = 8'h2d;    Blue = 8'h53;
end 12'he27:    begin Red = 8'h3e;    Green = 8'h23;    Blue = 8'h42;
end 12'he28:    begin Red = 8'h3b;    Green = 8'h1e;    Blue = 8'h3b;
end 12'he29:    begin Red = 8'h00;    Green = 8'h16;    Blue = 8'hf5;
end 12'he2a:    begin Red = 8'h4b;    Green = 8'h2b;    Blue = 8'h4d;
end 12'he2b:    begin Red = 8'h46;    Green = 8'h29;    Blue = 8'h46;
end 12'he2c:    begin Red = 8'hc7;    Green = 8'ha4;    Blue = 8'h56;
end 12'he2d:    begin Red = 8'h27;    Green = 8'h54;    Blue = 8'h72;
end 12'he2e:    begin Red = 8'h9a;    Green = 8'ha5;    Blue = 8'ha7;
end 12'he2f:    begin Red = 8'ha1;    Green = 8'ha4;    Blue = 8'ha6;
end 12'he30:    begin Red = 8'h80;    Green = 8'h89;    Blue = 8'h88;
end 12'he31:    begin Red = 8'h57;    Green = 8'hbe;    Blue = 8'hf2;
end 12'he32:    begin Red = 8'h55;    Green = 8'haf;    Blue = 8'hf4;
end 12'he33:    begin Red = 8'h18;    Green = 8'h5f;    Blue = 8'h95;
end 12'he34:    begin Red = 8'ha7;    Green = 8'hcb;    Blue = 8'h27;
end 12'he35:    begin Red = 8'he1;    Green = 8'he4;    Blue = 8'hd2;
end 12'he36:    begin Red = 8'h04;    Green = 8'h62;    Blue = 8'hd4;
end 12'he37:    begin Red = 8'h73;    Green = 8'h70;    Blue = 8'h3e;
end 12'he38:    begin Red = 8'h06;    Green = 8'h43;    Blue = 8'he8;
end 12'he39:    begin Red = 8'hae;    Green = 8'hd5;    Blue = 8'hd4;
end 12'he3a:    begin Red = 8'hbb;    Green = 8'h49;    Blue = 8'h38;
end 12'he3b:    begin Red = 8'hc4;    Green = 8'h61;    Blue = 8'h52;
end 12'he3c:    begin Red = 8'h48;    Green = 8'h30;    Blue = 8'h41;
end 12'he3d:    begin Red = 8'h42;    Green = 8'h2b;    Blue = 8'h39;
end 12'he3e:    begin Red = 8'hde;    Green = 8'hed;    Blue = 8'hac;
end 12'he3f:    begin Red = 8'h35;    Green = 8'h1c;    Blue = 8'h3a;
end 12'he40:    begin Red = 8'h39;    Green = 8'h1d;    Blue = 8'h41;
end 12'he41:    begin Red = 8'h01;    Green = 8'h01;    Blue = 8'h27;
end 12'he42:    begin Red = 8'h88;    Green = 8'h98;    Blue = 8'h9e;
end 12'he43:    begin Red = 8'h85;    Green = 8'h9d;    Blue = 8'h99;
end 12'he44:    begin Red = 8'h80;    Green = 8'h92;    Blue = 8'h9a;
end 12'he45:    begin Red = 8'h21;    Green = 8'h56;    Blue = 8'h98;
end 12'he46:    begin Red = 8'hb7;    Green = 8'hb6;    Blue = 8'h36;
end 12'he47:    begin Red = 8'hec;    Green = 8'hdc;    Blue = 8'hd7;
end 12'he48:    begin Red = 8'h88;    Green = 8'h81;    Blue = 8'h4b;
end 12'he49:    begin Red = 8'h78;    Green = 8'h76;    Blue = 8'h3f;
end 12'he4a:    begin Red = 8'h82;    Green = 8'h89;    Blue = 8'h95;
end 12'he4b:    begin Red = 8'h7d;    Green = 8'h95;    Blue = 8'h8f;
end 12'he4c:    begin Red = 8'hb8;    Green = 8'hd7;    Blue = 8'hc7;
end 12'he4d:    begin Red = 8'hb8;    Green = 8'hd4;    Blue = 8'hcd;
end 12'he4e:    begin Red = 8'hc5;    Green = 8'h44;    Blue = 8'h40;
end 12'he4f:    begin Red = 8'h51;    Green = 8'h2c;    Blue = 8'h55;
end 12'he50:    begin Red = 8'h41;    Green = 8'h24;    Blue = 8'h51;
end 12'he51:    begin Red = 8'h3f;    Green = 8'h23;    Blue = 8'h47;
end 12'he52:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'h06;
end 12'he53:    begin Red = 8'h45;    Green = 8'h29;    Blue = 8'h4e;
end 12'he54:    begin Red = 8'h3d;    Green = 8'h1f;    Blue = 8'h58;
end 12'he55:    begin Red = 8'h7a;    Green = 8'h65;    Blue = 8'h6d;
end 12'he56:    begin Red = 8'h72;    Green = 8'h5f;    Blue = 8'h68;
end 12'he57:    begin Red = 8'h47;    Green = 8'h2a;    Blue = 8'h55;
end 12'he58:    begin Red = 8'h36;    Green = 8'h1a;    Blue = 8'h4a;
end 12'he59:    begin Red = 8'h1b;    Green = 8'h1a;    Blue = 8'h17;
end 12'he5a:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'hd9;
end 12'he5b:    begin Red = 8'h55;    Green = 8'h48;    Blue = 8'h4a;
end 12'he5c:    begin Red = 8'h57;    Green = 8'h43;    Blue = 8'h48;
end 12'he5d:    begin Red = 8'h6a;    Green = 8'h92;    Blue = 8'h40;
end 12'he5e:    begin Red = 8'h69;    Green = 8'h8f;    Blue = 8'h46;
end 12'he5f:    begin Red = 8'h54;    Green = 8'h72;    Blue = 8'h38;
end 12'he60:    begin Red = 8'h38;    Green = 8'h5c;    Blue = 8'h19;
end 12'he61:    begin Red = 8'h8a;    Green = 8'h92;    Blue = 8'h98;
end 12'he62:    begin Red = 8'h10;    Green = 8'h1c;    Blue = 8'h29;
end 12'he63:    begin Red = 8'h1e;    Green = 8'h1c;    Blue = 8'h28;
end 12'he64:    begin Red = 8'h1c;    Green = 8'h20;    Blue = 8'h22;
end 12'he65:    begin Red = 8'h55;    Green = 8'h77;    Blue = 8'h86;
end 12'he66:    begin Red = 8'h54;    Green = 8'h32;    Blue = 8'h4b;
end 12'he67:    begin Red = 8'h22;    Green = 8'h16;    Blue = 8'h23;
end 12'he68:    begin Red = 8'h00;    Green = 8'h18;    Blue = 8'hfa;
end 12'he69:    begin Red = 8'h3b;    Green = 8'h2d;    Blue = 8'h38;
end 12'he6a:    begin Red = 8'h35;    Green = 8'h35;    Blue = 8'h25;
end 12'he6b:    begin Red = 8'h9e;    Green = 8'h97;    Blue = 8'h91;
end 12'he6c:    begin Red = 8'hb1;    Green = 8'hae;    Blue = 8'h99;
end 12'he6d:    begin Red = 8'h9e;    Green = 8'h92;    Blue = 8'h8e;
end 12'he6e:    begin Red = 8'h00;    Green = 8'h1d;    Blue = 8'h07;
end 12'he6f:    begin Red = 8'h02;    Green = 8'haa;    Blue = 8'h16;
end 12'he70:    begin Red = 8'h00;    Green = 8'h08;    Blue = 8'h00;
end 12'he71:    begin Red = 8'h00;    Green = 8'h08;    Blue = 8'h26;
end 12'he72:    begin Red = 8'h49;    Green = 8'h6f;    Blue = 8'h2b;
end 12'he73:    begin Red = 8'hf5;    Green = 8'he1;    Blue = 8'ha6;
end 12'he74:    begin Red = 8'he9;    Green = 8'hd2;    Blue = 8'h98;
end 12'he75:    begin Red = 8'h7c;    Green = 8'h73;    Blue = 8'h44;
end 12'he76:    begin Red = 8'h5c;    Green = 8'h53;    Blue = 8'h2d;
end 12'he77:    begin Red = 8'h63;    Green = 8'h33;    Blue = 8'h46;
end 12'he78:    begin Red = 8'h7a;    Green = 8'h76;    Blue = 8'h8f;
end 12'he79:    begin Red = 8'h01;    Green = 8'hf1;    Blue = 8'h0b;
end 12'he7a:    begin Red = 8'h3a;    Green = 8'h31;    Blue = 8'h3d;
end 12'he7b:    begin Red = 8'h02;    Green = 8'hcd;    Blue = 8'h1e;
end 12'he7c:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h2e;
end 12'he7d:    begin Red = 8'h1c;    Green = 8'h14;    Blue = 8'h10;
end 12'he7e:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h3e;
end 12'he7f:    begin Red = 8'h44;    Green = 8'h67;    Blue = 8'h27;
end 12'he80:    begin Red = 8'h64;    Green = 8'h69;    Blue = 8'h38;
end 12'he81:    begin Red = 8'h5c;    Green = 8'h63;    Blue = 8'h33;
end 12'he82:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'ha4;
end 12'he83:    begin Red = 8'h85;    Green = 8'h64;    Blue = 8'h17;
end 12'he84:    begin Red = 8'h2b;    Green = 8'h27;    Blue = 8'h33;
end 12'he85:    begin Red = 8'h08;    Green = 8'h35;    Blue = 8'hf4;
end 12'he86:    begin Red = 8'h56;    Green = 8'h3b;    Blue = 8'h3b;
end 12'he87:    begin Red = 8'hfd;    Green = 8'hf1;    Blue = 8'ha9;
end 12'he88:    begin Red = 8'h5b;    Green = 8'h2d;    Blue = 8'h65;
end 12'he89:    begin Red = 8'hc1;    Green = 8'hce;    Blue = 8'h90;
end 12'he8a:    begin Red = 8'h49;    Green = 8'h25;    Blue = 8'h5f;
end 12'he8b:    begin Red = 8'h55;    Green = 8'h2d;    Blue = 8'h65;
end 12'he8c:    begin Red = 8'h4f;    Green = 8'h27;    Blue = 8'h60;
end 12'he8d:    begin Red = 8'h00;    Green = 8'h1b;    Blue = 8'he5;
end 12'he8e:    begin Red = 8'h47;    Green = 8'h24;    Blue = 8'h57;
end 12'he8f:    begin Red = 8'h50;    Green = 8'h23;    Blue = 8'h5b;
end 12'he90:    begin Red = 8'h41;    Green = 8'h7a;    Blue = 8'h3f;
end 12'he91:    begin Red = 8'h6c;    Green = 8'h66;    Blue = 8'h5e;
end 12'he92:    begin Red = 8'h5e;    Green = 8'h3d;    Blue = 8'h24;
end 12'he93:    begin Red = 8'h02;    Green = 8'h87;    Blue = 8'h19;
end 12'he94:    begin Red = 8'h01;    Green = 8'h31;    Blue = 8'h2d;
end 12'he95:    begin Red = 8'h01;    Green = 8'h21;    Blue = 8'h1e;
end 12'he96:    begin Red = 8'h01;    Green = 8'ha1;    Blue = 8'h2e;
end 12'he97:    begin Red = 8'h01;    Green = 8'hb1;    Blue = 8'h1e;
end 12'he98:    begin Red = 8'h56;    Green = 8'h76;    Blue = 8'h30;
end 12'he99:    begin Red = 8'he3;    Green = 8'hcf;    Blue = 8'h9c;
end 12'he9a:    begin Red = 8'h8a;    Green = 8'h88;    Blue = 8'h4b;
end 12'he9b:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'hc4;
end 12'he9c:    begin Red = 8'h33;    Green = 8'h2e;    Blue = 8'h3b;
end 12'he9d:    begin Red = 8'h07;    Green = 8'hf5;    Blue = 8'hfe;
end 12'he9e:    begin Red = 8'h08;    Green = 8'h25;    Blue = 8'hf6;
end 12'he9f:    begin Red = 8'hb9;    Green = 8'hc9;    Blue = 8'h88;
end 12'hea0:    begin Red = 8'h38;    Green = 8'h21;    Blue = 8'h6d;
end 12'hea1:    begin Red = 8'h33;    Green = 8'h22;    Blue = 8'h6c;
end 12'hea2:    begin Red = 8'h2d;    Green = 8'h1c;    Blue = 8'h66;
end 12'hea3:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h55;
end 12'hea4:    begin Red = 8'h3a;    Green = 8'h8c;    Blue = 8'h3e;
end 12'hea5:    begin Red = 8'h00;    Green = 8'h20;    Blue = 8'h0e;
end 12'hea6:    begin Red = 8'h00;    Green = 8'h09;    Blue = 8'h56;
end 12'hea7:    begin Red = 8'h01;    Green = 8'h51;    Blue = 8'h2d;
end 12'hea8:    begin Red = 8'h17;    Green = 8'h11;    Blue = 8'h12;
end 12'hea9:    begin Red = 8'h00;    Green = 8'h0a;    Blue = 8'h05;
end 12'heaa:    begin Red = 8'h98;    Green = 8'had;    Blue = 8'ha1;
end 12'heab:    begin Red = 8'h04;    Green = 8'he2;    Blue = 8'he3;
end 12'heac:    begin Red = 8'h04;    Green = 8'h42;    Blue = 8'hd4;
end 12'head:    begin Red = 8'h92;    Green = 8'ha5;    Blue = 8'ha6;
end 12'heae:    begin Red = 8'h74;    Green = 8'h76;    Blue = 8'h81;
end 12'heaf:    begin Red = 8'h5c;    Green = 8'h41;    Blue = 8'h41;
end 12'heb0:    begin Red = 8'h5c;    Green = 8'h39;    Blue = 8'h4f;
end 12'heb1:    begin Red = 8'hc1;    Green = 8'ha9;    Blue = 8'h6e;
end 12'heb2:    begin Red = 8'h5e;    Green = 8'h2d;    Blue = 8'h6b;
end 12'heb3:    begin Red = 8'h50;    Green = 8'h27;    Blue = 8'h65;
end 12'heb4:    begin Red = 8'h58;    Green = 8'h2d;    Blue = 8'h6a;
end 12'heb5:    begin Red = 8'h00;    Green = 8'h19;    Blue = 8'hd1;
end 12'heb6:    begin Red = 8'h4f;    Green = 8'h2d;    Blue = 8'h64;
end 12'heb7:    begin Red = 8'hc0;    Green = 8'h3d;    Blue = 8'h2f;
end 12'heb8:    begin Red = 8'h49;    Green = 8'h29;    Blue = 8'h66;
end 12'heb9:    begin Red = 8'h00;    Green = 8'he8;    Blue = 8'h22;
end 12'heba:    begin Red = 8'h00;    Green = 8'hdd;    Blue = 8'ha3;
end 12'hebb:    begin Red = 8'h2a;    Green = 8'h19;    Blue = 8'h10;
end 12'hebc:    begin Red = 8'h50;    Green = 8'h7c;    Blue = 8'h36;
end 12'hebd:    begin Red = 8'h51;    Green = 8'h74;    Blue = 8'h33;
end 12'hebe:    begin Red = 8'h39;    Green = 8'h86;    Blue = 8'h47;
end 12'hebf:    begin Red = 8'h87;    Green = 8'hb0;    Blue = 8'ha5;
end 12'hec0:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'hc0;
end 12'hec1:    begin Red = 8'h0b;    Green = 8'hf2;    Blue = 8'h7e;
end 12'hec2:    begin Red = 8'hb3;    Green = 8'h27;    Blue = 8'h17;
end 12'hec3:    begin Red = 8'hba;    Green = 8'h2c;    Blue = 8'h15;
end 12'hec4:    begin Red = 8'hbf;    Green = 8'h28;    Blue = 8'h20;
end 12'hec5:    begin Red = 8'hc3;    Green = 8'h25;    Blue = 8'h19;
end 12'hec6:    begin Red = 8'hb8;    Green = 8'h25;    Blue = 8'h1a;
end 12'hec7:    begin Red = 8'hb9;    Green = 8'h23;    Blue = 8'h21;
end 12'hec8:    begin Red = 8'h8d;    Green = 8'h21;    Blue = 8'h14;
end 12'hec9:    begin Red = 8'h88;    Green = 8'h19;    Blue = 8'h11;
end 12'heca:    begin Red = 8'h82;    Green = 8'h23;    Blue = 8'h10;
end 12'hecb:    begin Red = 8'h5f;    Green = 8'h4b;    Blue = 8'h64;
end 12'hecc:    begin Red = 8'h56;    Green = 8'h4b;    Blue = 8'h62;
end 12'hecd:    begin Red = 8'h46;    Green = 8'h1f;    Blue = 8'h5d;
end 12'hece:    begin Red = 8'h38;    Green = 8'h1b;    Blue = 8'h5b;
end 12'hecf:    begin Red = 8'h2c;    Green = 8'h1c;    Blue = 8'h5a;
end 12'hed0:    begin Red = 8'h5b;    Green = 8'h27;    Blue = 8'h6b;
end 12'hed1:    begin Red = 8'h32;    Green = 8'h18;    Blue = 8'h54;
end 12'hed2:    begin Red = 8'h58;    Green = 8'h24;    Blue = 8'h73;
end 12'hed3:    begin Red = 8'h37;    Green = 8'h17;    Blue = 8'h55;
end 12'hed4:    begin Red = 8'h00;    Green = 8'hf2;    Blue = 8'h46;
end 12'hed5:    begin Red = 8'h1c;    Green = 8'h5a;    Blue = 8'h82;
end 12'hed6:    begin Red = 8'h21;    Green = 8'h5c;    Blue = 8'h96;
end 12'hed7:    begin Red = 8'h27;    Green = 8'h4e;    Blue = 8'h7c;
end 12'hed8:    begin Red = 8'h9b;    Green = 8'h88;    Blue = 8'h8f;
end 12'hed9:    begin Red = 8'h00;    Green = 8'hea;    Blue = 8'h03;
end 12'heda:    begin Red = 8'h00;    Green = 8'he1;    Blue = 8'h6e;
end 12'hedb:    begin Red = 8'h68;    Green = 8'h9b;    Blue = 8'h41;
end 12'hedc:    begin Red = 8'h65;    Green = 8'h45;    Blue = 8'h3f;
end 12'hedd:    begin Red = 8'h73;    Green = 8'h5c;    Blue = 8'h44;
end 12'hede:    begin Red = 8'h53;    Green = 8'h72;    Blue = 8'h3f;
end 12'hedf:    begin Red = 8'h4c;    Green = 8'h69;    Blue = 8'h32;
end 12'hee0:    begin Red = 8'h32;    Green = 8'h88;    Blue = 8'h4a;
end 12'hee1:    begin Red = 8'h00;    Green = 8'he4;    Blue = 8'hb6;
end 12'hee2:    begin Red = 8'h87;    Green = 8'hae;    Blue = 8'h9d;
end 12'hee3:    begin Red = 8'hcc;    Green = 8'hbd;    Blue = 8'h8d;
end 12'hee4:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'h61;
end 12'hee5:    begin Red = 8'h04;    Green = 8'h62;    Blue = 8'h97;
end 12'hee6:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h57;
end 12'hee7:    begin Red = 8'h3e;    Green = 8'h3c;    Blue = 8'h43;
end 12'hee8:    begin Red = 8'h0c;    Green = 8'h3d;    Blue = 8'h43;
end 12'hee9:    begin Red = 8'hba;    Green = 8'h2b;    Blue = 8'h1c;
end 12'heea:    begin Red = 8'hbd;    Green = 8'h27;    Blue = 8'h15;
end 12'heeb:    begin Red = 8'h83;    Green = 8'h21;    Blue = 8'h17;
end 12'heec:    begin Red = 8'he3;    Green = 8'hcf;    Blue = 8'ha3;
end 12'heed:    begin Red = 8'he7;    Green = 8'hf2;    Blue = 8'hb4;
end 12'heee:    begin Red = 8'h34;    Green = 8'h1a;    Blue = 8'h60;
end 12'heef:    begin Red = 8'h33;    Green = 8'h1d;    Blue = 8'h5a;
end 12'hef0:    begin Red = 8'h4f;    Green = 8'h2e;    Blue = 8'h6a;
end 12'hef1:    begin Red = 8'hc0;    Green = 8'h3e;    Blue = 8'h38;
end 12'hef2:    begin Red = 8'hb8;    Green = 8'h3e;    Blue = 8'h2b;
end 12'hef3:    begin Red = 8'h58;    Green = 8'h2d;    Blue = 8'h60;
end 12'hef4:    begin Red = 8'h6d;    Green = 8'h60;    Blue = 8'h5e;
end 12'hef5:    begin Red = 8'h20;    Green = 8'h52;    Blue = 8'h7e;
end 12'hef6:    begin Red = 8'h98;    Green = 8'h93;    Blue = 8'h81;
end 12'hef7:    begin Red = 8'h00;    Green = 8'hf3;    Blue = 8'h03;
end 12'hef8:    begin Red = 8'h70;    Green = 8'h8c;    Blue = 8'h46;
end 12'hef9:    begin Red = 8'h70;    Green = 8'ha0;    Blue = 8'h5a;
end 12'hefa:    begin Red = 8'h2f;    Green = 8'h87;    Blue = 8'h41;
end 12'hefb:    begin Red = 8'h0d;    Green = 8'ha8;    Blue = 8'h12;
end 12'hefc:    begin Red = 8'h8e;    Green = 8'hb4;    Blue = 8'ha8;
end 12'hefd:    begin Red = 8'h02;    Green = 8'he1;    Blue = 8'h45;
end 12'hefe:    begin Red = 8'h06;    Green = 8'hb4;    Blue = 8'h1c;
end 12'heff:    begin Red = 8'hd6;    Green = 8'ha9;    Blue = 8'h84;
end 12'hf00:    begin Red = 8'h74;    Green = 8'h81;    Blue = 8'h5e;
end 12'hf01:    begin Red = 8'h52;    Green = 8'h54;    Blue = 8'h72;
end 12'hf02:    begin Red = 8'h4e;    Green = 8'h4e;    Blue = 8'h77;
end 12'hf03:    begin Red = 8'h33;    Green = 8'h30;    Blue = 8'h47;
end 12'hf04:    begin Red = 8'h16;    Green = 8'h32;    Blue = 8'h50;
end 12'hf05:    begin Red = 8'h0b;    Green = 8'h22;    Blue = 8'haf;
end 12'hf06:    begin Red = 8'h8e;    Green = 8'h1b;    Blue = 8'h13;
end 12'hf07:    begin Red = 8'h60;    Green = 8'h50;    Blue = 8'h63;
end 12'hf08:    begin Red = 8'h62;    Green = 8'h43;    Blue = 8'h44;
end 12'hf09:    begin Red = 8'h63;    Green = 8'h41;    Blue = 8'h50;
end 12'hf0a:    begin Red = 8'hea;    Green = 8'hf2;    Blue = 8'hc3;
end 12'hf0b:    begin Red = 8'hbb;    Green = 8'h3e;    Blue = 8'h31;
end 12'hf0c:    begin Red = 8'h15;    Green = 8'h4d;    Blue = 8'h8e;
end 12'hf0d:    begin Red = 8'h07;    Green = 8'h48;    Blue = 8'h81;
end 12'hf0e:    begin Red = 8'h3e;    Green = 8'h59;    Blue = 8'h1f;
end 12'hf0f:    begin Red = 8'h4c;    Green = 8'h63;    Blue = 8'h32;
end 12'hf10:    begin Red = 8'h7b;    Green = 8'hab;    Blue = 8'h53;
end 12'hf11:    begin Red = 8'h52;    Green = 8'hba;    Blue = 8'he8;
end 12'hf12:    begin Red = 8'hd6;    Green = 8'haf;    Blue = 8'h79;
end 12'hf13:    begin Red = 8'hdc;    Green = 8'hb5;    Blue = 8'h7e;
end 12'hf14:    begin Red = 8'h05;    Green = 8'h33;    Blue = 8'h24;
end 12'hf15:    begin Red = 8'hef;    Green = 8'hef;    Blue = 8'hbe;
end 12'hf16:    begin Red = 8'h6a;    Green = 8'h89;    Blue = 8'h59;
end 12'hf17:    begin Red = 8'h0d;    Green = 8'h01;    Blue = 8'h5c;
end 12'hf18:    begin Red = 8'h57;    Green = 8'h4b;    Blue = 8'h73;
end 12'hf19:    begin Red = 8'h44;    Green = 8'h4a;    Blue = 8'h75;
end 12'hf1a:    begin Red = 8'h50;    Green = 8'h4f;    Blue = 8'h64;
end 12'hf1b:    begin Red = 8'h5c;    Green = 8'h5a;    Blue = 8'h79;
end 12'hf1c:    begin Red = 8'hb1;    Green = 8'h24;    Blue = 8'h11;
end 12'hf1d:    begin Red = 8'hb3;    Green = 8'h2d;    Blue = 8'h1c;
end 12'hf1e:    begin Red = 8'h08;    Green = 8'h31;    Blue = 8'h99;
end 12'hf1f:    begin Red = 8'h76;    Green = 8'h1e;    Blue = 8'h1b;
end 12'hf20:    begin Red = 8'h5d;    Green = 8'h57;    Blue = 8'h74;
end 12'hf21:    begin Red = 8'h56;    Green = 8'h59;    Blue = 8'h7b;
end 12'hf22:    begin Red = 8'h58;    Green = 8'h50;    Blue = 8'h79;
end 12'hf23:    begin Red = 8'h00;    Green = 8'h07;    Blue = 8'h32;
end 12'hf24:    begin Red = 8'hbc;    Green = 8'h26;    Blue = 8'h26;
end 12'hf25:    begin Red = 8'hc4;    Green = 8'h30;    Blue = 8'h26;
end 12'hf26:    begin Red = 8'hd4;    Green = 8'h3e;    Blue = 8'h36;
end 12'hf27:    begin Red = 8'hba;    Green = 8'h2a;    Blue = 8'h21;
end 12'hf28:    begin Red = 8'haa;    Green = 8'h2b;    Blue = 8'h21;
end 12'hf29:    begin Red = 8'h4f;    Green = 8'h52;    Blue = 8'h43;
end 12'hf2a:    begin Red = 8'h26;    Green = 8'h53;    Blue = 8'h8d;
end 12'hf2b:    begin Red = 8'h00;    Green = 8'h27;    Blue = 8'h90;
end 12'hf2c:    begin Red = 8'h00;    Green = 8'h29;    Blue = 8'h00;
end 12'hf2d:    begin Red = 8'h1d;    Green = 8'h55;    Blue = 8'h86;
end 12'hf2e:    begin Red = 8'ha0;    Green = 8'h89;    Blue = 8'h8d;
end 12'hf2f:    begin Red = 8'h78;    Green = 8'h6b;    Blue = 8'h74;
end 12'hf30:    begin Red = 8'h74;    Green = 8'h65;    Blue = 8'h71;
end 12'hf31:    begin Red = 8'h73;    Green = 8'h65;    Blue = 8'h6b;
end 12'hf32:    begin Red = 8'hd3;    Green = 8'hc5;    Blue = 8'h92;
end 12'hf33:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'h25;
end 12'hf34:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'h88;
end 12'hf35:    begin Red = 8'hc2;    Green = 8'ha2;    Blue = 8'h6a;
end 12'hf36:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h83;
end 12'hf37:    begin Red = 8'he3;    Green = 8'he6;    Blue = 8'hb7;
end 12'hf38:    begin Red = 8'h0d;    Green = 8'h01;    Blue = 8'hc3;
end 12'hf39:    begin Red = 8'h83;    Green = 8'h1a;    Blue = 8'h16;
end 12'hf3a:    begin Red = 8'h87;    Green = 8'h20;    Blue = 8'h10;
end 12'hf3b:    begin Red = 8'h40;    Green = 8'h2b;    Blue = 8'h60;
end 12'hf3c:    begin Red = 8'hb0;    Green = 8'h9d;    Blue = 8'h64;
end 12'hf3d:    begin Red = 8'h0d;    Green = 8'h44;    Blue = 8'h7e;
end 12'hf3e:    begin Red = 8'hff;    Green = 8'hfa;    Blue = 8'hf0;
end 12'hf3f:    begin Red = 8'h00;    Green = 8'h30;    Blue = 8'h6b;
end 12'hf40:    begin Red = 8'h21;    Green = 8'h51;    Blue = 8'h77;
end 12'hf41:    begin Red = 8'h1e;    Green = 8'h6d;    Blue = 8'had;
end 12'hf42:    begin Red = 8'h25;    Green = 8'h69;    Blue = 8'haf;
end 12'hf43:    begin Red = 8'h25;    Green = 8'h69;    Blue = 8'ha7;
end 12'hf44:    begin Red = 8'h28;    Green = 8'hfa;    Blue = 8'hf6;
end 12'hf45:    begin Red = 8'h25;    Green = 8'hf3;    Blue = 8'hf2;
end 12'hf46:    begin Red = 8'h24;    Green = 8'h2e;    Blue = 8'h6d;
end 12'hf47:    begin Red = 8'h23;    Green = 8'h56;    Blue = 8'h84;
end 12'hf48:    begin Red = 8'h13;    Green = 8'h3e;    Blue = 8'h68;
end 12'hf49:    begin Red = 8'h3e;    Green = 8'h59;    Blue = 8'h2f;
end 12'hf4a:    begin Red = 8'hc8;    Green = 8'h97;    Blue = 8'h62;
end 12'hf4b:    begin Red = 8'h7e;    Green = 8'h71;    Blue = 8'h55;
end 12'hf4c:    begin Red = 8'hb5;    Green = 8'h2d;    Blue = 8'h16;
end 12'hf4d:    begin Red = 8'h94;    Green = 8'h20;    Blue = 8'h12;
end 12'hf4e:    begin Red = 8'ha0;    Green = 8'h20;    Blue = 8'h12;
end 12'hf4f:    begin Red = 8'h96;    Green = 8'h1f;    Blue = 8'h1a;
end 12'hf50:    begin Red = 8'h99;    Green = 8'h1f;    Blue = 8'h11;
end 12'hf51:    begin Red = 8'hff;    Green = 8'h8f;    Blue = 8'h1c;
end 12'hf52:    begin Red = 8'hfb;    Green = 8'h78;    Blue = 8'h24;
end 12'hf53:    begin Red = 8'hfe;    Green = 8'h80;    Blue = 8'h23;
end 12'hf54:    begin Red = 8'hf6;    Green = 8'h7d;    Blue = 8'h1e;
end 12'hf55:    begin Red = 8'haa;    Green = 8'h9c;    Blue = 8'h68;
end 12'hf56:    begin Red = 8'h44;    Green = 8'h25;    Blue = 8'h22;
end 12'hf57:    begin Red = 8'h1f;    Green = 8'h69;    Blue = 8'ha7;
end 12'hf58:    begin Red = 8'h23;    Green = 8'h70;    Blue = 8'hab;
end 12'hf59:    begin Red = 8'h25;    Green = 8'h64;    Blue = 8'hb6;
end 12'hf5a:    begin Red = 8'h30;    Green = 8'hf4;    Blue = 8'hf5;
end 12'hf5b:    begin Red = 8'h1f;    Green = 8'hfa;    Blue = 8'hf6;
end 12'hf5c:    begin Red = 8'h24;    Green = 8'h5c;    Blue = 8'h85;
end 12'hf5d:    begin Red = 8'h23;    Green = 8'hf3;    Blue = 8'he8;
end 12'hf5e:    begin Red = 8'h8d;    Green = 8'h85;    Blue = 8'h7a;
end 12'hf5f:    begin Red = 8'h45;    Green = 8'h59;    Blue = 8'h2f;
end 12'hf60:    begin Red = 8'h72;    Green = 8'h92;    Blue = 8'h46;
end 12'hf61:    begin Red = 8'h6f;    Green = 8'h90;    Blue = 8'h4f;
end 12'hf62:    begin Red = 8'h51;    Green = 8'h6f;    Blue = 8'h33;
end 12'hf63:    begin Red = 8'h4c;    Green = 8'h65;    Blue = 8'h37;
end 12'hf64:    begin Red = 8'h5f;    Green = 8'h75;    Blue = 8'h3e;
end 12'hf65:    begin Red = 8'h63;    Green = 8'h6a;    Blue = 8'h30;
end 12'hf66:    begin Red = 8'h6d;    Green = 8'h6a;    Blue = 8'h36;
end 12'hf67:    begin Red = 8'hce;    Green = 8'h28;    Blue = 8'h19;
end 12'hf68:    begin Red = 8'hd4;    Green = 8'h28;    Blue = 8'h13;
end 12'hf69:    begin Red = 8'h00;    Green = 8'hd5;    Blue = 8'h20;
end 12'hf6a:    begin Red = 8'ha0;    Green = 8'h1c;    Blue = 8'h19;
end 12'hf6b:    begin Red = 8'h09;    Green = 8'h12;    Blue = 8'h1d;
end 12'hf6c:    begin Red = 8'h0b;    Green = 8'hb2;    Blue = 8'hab;
end 12'hf6d:    begin Red = 8'hcd;    Green = 8'h24;    Blue = 8'h10;
end 12'hf6e:    begin Red = 8'hda;    Green = 8'h28;    Blue = 8'h19;
end 12'hf6f:    begin Red = 8'h0b;    Green = 8'he1;    Blue = 8'h10;
end 12'hf70:    begin Red = 8'h00;    Green = 8'hd4;    Blue = 8'h00;
end 12'hf71:    begin Red = 8'hfb;    Green = 8'ha3;    Blue = 8'h2c;
end 12'hf72:    begin Red = 8'h45;    Green = 8'h23;    Blue = 8'h39;
end 12'hf73:    begin Red = 8'h4c;    Green = 8'h4b;    Blue = 8'h51;
end 12'hf74:    begin Red = 8'h3d;    Green = 8'h23;    Blue = 8'h21;
end 12'hf75:    begin Red = 8'h21;    Green = 8'h6b;    Blue = 8'hb7;
end 12'hf76:    begin Red = 8'h24;    Green = 8'h64;    Blue = 8'haf;
end 12'hf77:    begin Red = 8'h22;    Green = 8'h5f;    Blue = 8'haf;
end 12'hf78:    begin Red = 8'h1b;    Green = 8'h49;    Blue = 8'h9d;
end 12'hf79:    begin Red = 8'h1d;    Green = 8'hf9;    Blue = 8'hf1;
end 12'hf7a:    begin Red = 8'h1f;    Green = 8'hee;    Blue = 8'hdc;
end 12'hf7b:    begin Red = 8'h46;    Green = 8'h6e;    Blue = 8'h35;
end 12'hf7c:    begin Red = 8'h75;    Green = 8'ha3;    Blue = 8'h4e;
end 12'hf7d:    begin Red = 8'h6f;    Green = 8'hac;    Blue = 8'h50;
end 12'hf7e:    begin Red = 8'h55;    Green = 8'h7f;    Blue = 8'h36;
end 12'hf7f:    begin Red = 8'h55;    Green = 8'h82;    Blue = 8'h41;
end 12'hf80:    begin Red = 8'h05;    Green = 8'h02;    Blue = 8'h84;
end 12'hf81:    begin Red = 8'h76;    Green = 8'h84;    Blue = 8'h4b;
end 12'hf82:    begin Red = 8'h52;    Green = 8'h63;    Blue = 8'h30;
end 12'hf83:    begin Red = 8'h06;    Green = 8'hb3;    Blue = 8'h92;
end 12'hf84:    begin Red = 8'h62;    Green = 8'h6c;    Blue = 8'h43;
end 12'hf85:    begin Red = 8'h40;    Green = 8'h57;    Blue = 8'h25;
end 12'hf86:    begin Red = 8'hb8;    Green = 8'h25;    Blue = 8'h12;
end 12'hf87:    begin Red = 8'hbf;    Green = 8'h2c;    Blue = 8'h17;
end 12'hf88:    begin Red = 8'h0f;    Green = 8'h15;    Blue = 8'h12;
end 12'hf89:    begin Red = 8'h25;    Green = 8'heb;    Blue = 8'hf0;
end 12'hf8a:    begin Red = 8'h40;    Green = 8'hdb;    Blue = 8'hf6;
end 12'hf8b:    begin Red = 8'h9d;    Green = 8'h77;    Blue = 8'h63;
end 12'hf8c:    begin Red = 8'h07;    Green = 8'hb1;    Blue = 8'hee;
end 12'hf8d:    begin Red = 8'h1d;    Green = 8'h53;    Blue = 8'h9e;
end 12'hf8e:    begin Red = 8'h30;    Green = 8'hef;    Blue = 8'hf3;
end 12'hf8f:    begin Red = 8'h26;    Green = 8'hf5;    Blue = 8'hed;
end 12'hf90:    begin Red = 8'h48;    Green = 8'h3c;    Blue = 8'h1c;
end 12'hf91:    begin Red = 8'h46;    Green = 8'h28;    Blue = 8'h1c;
end 12'hf92:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'hc5;
end 12'hf93:    begin Red = 8'h07;    Green = 8'h24;    Blue = 8'h39;
end 12'hf94:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'hd6;
end 12'hf95:    begin Red = 8'h04;    Green = 8'h42;    Blue = 8'h59;
end 12'hf96:    begin Red = 8'h05;    Green = 8'h93;    Blue = 8'h26;
end 12'hf97:    begin Red = 8'h08;    Green = 8'h81;    Blue = 8'h8d;
end 12'hf98:    begin Red = 8'ha4;    Green = 8'h79;    Blue = 8'h61;
end 12'hf99:    begin Red = 8'h7c;    Green = 8'h23;    Blue = 8'h10;
end 12'hf9a:    begin Red = 8'h7b;    Green = 8'h1d;    Blue = 8'h12;
end 12'hf9b:    begin Red = 8'h09;    Green = 8'h41;    Blue = 8'hae;
end 12'hf9c:    begin Red = 8'h05;    Green = 8'h15;    Blue = 8'h14;
end 12'hf9d:    begin Red = 8'h48;    Green = 8'h1d;    Blue = 8'h36;
end 12'hf9e:    begin Red = 8'h00;    Green = 8'hc5;    Blue = 8'h14;
end 12'hf9f:    begin Red = 8'h03;    Green = 8'hc2;    Blue = 8'h56;
end 12'hfa0:    begin Red = 8'h24;    Green = 8'h59;    Blue = 8'h7c;
end 12'hfa1:    begin Red = 8'h00;    Green = 8'h0d;    Blue = 8'h0a;
end 12'hfa2:    begin Red = 8'h1d;    Green = 8'h2f;    Blue = 8'h67;
end 12'hfa3:    begin Red = 8'h44;    Green = 8'h2a;    Blue = 8'h12;
end 12'hfa4:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'ha0;
end 12'hfa5:    begin Red = 8'hbe;    Green = 8'had;    Blue = 8'h83;
end 12'hfa6:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h70;
end 12'hfa7:    begin Red = 8'h03;    Green = 8'h91;    Blue = 8'he1;
end 12'hfa8:    begin Red = 8'h03;    Green = 8'ha1;    Blue = 8'hf1;
end 12'hfa9:    begin Red = 8'h02;    Green = 8'h41;    Blue = 8'h52;
end 12'hfaa:    begin Red = 8'h03;    Green = 8'h31;    Blue = 8'h90;
end 12'hfab:    begin Red = 8'h08;    Green = 8'h81;    Blue = 8'hcf;
end 12'hfac:    begin Red = 8'h14;    Green = 8'h15;    Blue = 8'h19;
end 12'hfad:    begin Red = 8'h99;    Green = 8'h26;    Blue = 8'h13;
end 12'hfae:    begin Red = 8'h31;    Green = 8'h15;    Blue = 8'h11;
end 12'hfaf:    begin Red = 8'h00;    Green = 8'h0a;    Blue = 8'h20;
end 12'hfb0:    begin Red = 8'h1c;    Green = 8'h11;    Blue = 8'h1e;
end 12'hfb1:    begin Red = 8'h10;    Green = 8'h12;    Blue = 8'h26;
end 12'hfb2:    begin Red = 8'h10;    Green = 8'h14;    Blue = 8'h2d;
end 12'hfb3:    begin Red = 8'h01;    Green = 8'h6d;    Blue = 8'h29;
end 12'hfb4:    begin Red = 8'h21;    Green = 8'h52;    Blue = 8'h8b;
end 12'hfb5:    begin Red = 8'h02;    Green = 8'hf1;    Blue = 8'hb3;
end 12'hfb6:    begin Red = 8'hf3;    Green = 8'hbf;    Blue = 8'h80;
end 12'hfb7:    begin Red = 8'h02;    Green = 8'h91;    Blue = 8'h84;
end 12'hfb8:    begin Red = 8'h00;    Green = 8'h15;    Blue = 8'h12;
end 12'hfb9:    begin Red = 8'h03;    Green = 8'h61;    Blue = 8'hf0;
end 12'hfba:    begin Red = 8'h03;    Green = 8'h72;    Blue = 8'h01;
end 12'hfbb:    begin Red = 8'h43;    Green = 8'hb1;    Blue = 8'hf3;
end 12'hfbc:    begin Red = 8'h43;    Green = 8'h98;    Blue = 8'he2;
end 12'hfbd:    begin Red = 8'h38;    Green = 8'h95;    Blue = 8'he3;
end 12'hfbe:    begin Red = 8'hc6;    Green = 8'hc1;    Blue = 8'h8b;
end 12'hfbf:    begin Red = 8'hd9;    Green = 8'hcc;    Blue = 8'h9c;
end 12'hfc0:    begin Red = 8'h1a;    Green = 8'h19;    Blue = 8'h36;
end 12'hfc1:    begin Red = 8'h0b;    Green = 8'h16;    Blue = 8'h32;
end 12'hfc2:    begin Red = 8'h1b;    Green = 8'h20;    Blue = 8'h1b;
end 12'hfc3:    begin Red = 8'hac;    Green = 8'hf4;    Blue = 8'hf4;
end 12'hfc4:    begin Red = 8'h00;    Green = 8'h00;    Blue = 8'h20;
end 12'hfc5:    begin Red = 8'hc4;    Green = 8'hf6;    Blue = 8'hf4;
end 12'hfc6:    begin Red = 8'ha0;    Green = 8'hfc;    Blue = 8'hf5;
end 12'hfc7:    begin Red = 8'h4c;    Green = 8'h4d;    Blue = 8'h58;
end 12'hfc8:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'hb5;
end 12'hfc9:    begin Red = 8'hfa;    Green = 8'hbd;    Blue = 8'h75;
end 12'hfca:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'ha1;
end 12'hfcb:    begin Red = 8'h03;    Green = 8'h81;    Blue = 8'hd0;
end 12'hfcc:    begin Red = 8'h4c;    Green = 8'h34;    Blue = 8'h12;
end 12'hfcd:    begin Red = 8'h3a;    Green = 8'hbe;    Blue = 8'hf6;
end 12'hfce:    begin Red = 8'h3a;    Green = 8'hb4;    Blue = 8'hf4;
end 12'hfcf:    begin Red = 8'h3d;    Green = 8'hc3;    Blue = 8'hf6;
end 12'hfd0:    begin Red = 8'h02;    Green = 8'h82;    Blue = 8'h15;
end 12'hfd1:    begin Red = 8'h97;    Green = 8'h83;    Blue = 8'h56;
end 12'hfd2:    begin Red = 8'h49;    Green = 8'h4e;    Blue = 8'h43;
end 12'hfd3:    begin Red = 8'h6b;    Green = 8'h5c;    Blue = 8'h66;
end 12'hfd4:    begin Red = 8'hc9;    Green = 8'hfc;    Blue = 8'hf5;
end 12'hfd5:    begin Red = 8'h57;    Green = 8'h50;    Blue = 8'h52;
end 12'hfd6:    begin Red = 8'h55;    Green = 8'h49;    Blue = 8'h4f;
end 12'hfd7:    begin Red = 8'hc4;    Green = 8'hfb;    Blue = 8'hf6;
end 12'hfd8:    begin Red = 8'h3c;    Green = 8'h46;    Blue = 8'h3d;
end 12'hfd9:    begin Red = 8'h3a;    Green = 8'hab;    Blue = 8'hf6;
end 12'hfda:    begin Red = 8'h37;    Green = 8'h96;    Blue = 8'hdd;
end 12'hfdb:    begin Red = 8'h33;    Green = 8'haa;    Blue = 8'hf5;
end 12'hfdc:    begin Red = 8'h67;    Green = 8'h63;    Blue = 8'h5c;
end 12'hfdd:    begin Red = 8'h6b;    Green = 8'h5a;    Blue = 8'h5b;
end 12'hfde:    begin Red = 8'hb6;    Green = 8'hfc;    Blue = 8'hf7;
end 12'hfdf:    begin Red = 8'ha7;    Green = 8'hfc;    Blue = 8'hf7;
end 12'hfe0:    begin Red = 8'h63;    Green = 8'h66;    Blue = 8'h53;
end 12'hfe1:    begin Red = 8'h6b;    Green = 8'h69;    Blue = 8'h64;
end 12'hfe2:    begin Red = 8'h5d;    Green = 8'h5c;    Blue = 8'h66;
end 12'hfe3:    begin Red = 8'h6a;    Green = 8'h60;    Blue = 8'h57;
end 12'hfe4:    begin Red = 8'h63;    Green = 8'h57;    Blue = 8'h66;
end 12'hfe5:    begin Red = 8'h62;    Green = 8'h60;    Blue = 8'h66;
end 12'hfe6:    begin Red = 8'h61;    Green = 8'h63;    Blue = 8'h71;
end 12'hfe7:    begin Red = 8'h5d;    Green = 8'h63;    Blue = 8'h69;
end 12'hfe8:    begin Red = 8'h6c;    Green = 8'h5e;    Blue = 8'h6d;
end 12'hfe9:    begin Red = 8'h5c;    Green = 8'h62;    Blue = 8'h6f;
end 12'hfea:    begin Red = 8'h54;    Green = 8'h62;    Blue = 8'h63;
end 12'hfeb:    begin Red = 8'h9e;    Green = 8'h86;    Blue = 8'h35;
end 12'hfec:    begin Red = 8'ha9;    Green = 8'h8f;    Blue = 8'h24;
end 12'hfed:    begin Red = 8'h70;    Green = 8'h70;    Blue = 8'h5c;
end 12'hfee:    begin Red = 8'ha0;    Green = 8'h82;    Blue = 8'h26;
end 12'hfef:    begin Red = 8'ha3;    Green = 8'h87;    Blue = 8'h29;
end 12'hff0:    begin Red = 8'h76;    Green = 8'h70;    Blue = 8'h68;
end 12'hff1:    begin Red = 8'hbe;    Green = 8'hc4;    Blue = 8'h92;
end 12'hff2:    begin Red = 8'h71;    Green = 8'h71;    Blue = 8'h61;
end 12'hff3:    begin Red = 8'hcd;    Green = 8'hb8;    Blue = 8'h98;
end 12'hff4:    begin Red = 8'hbf;    Green = 8'hae;    Blue = 8'h88;
end 12'hff5:    begin Red = 8'hb5;    Green = 8'ha4;    Blue = 8'h7e;
end 12'hff6:    begin Red = 8'haf;    Green = 8'h9f;    Blue = 8'h7c;
end 12'hff7:    begin Red = 8'had;    Green = 8'h9b;    Blue = 8'h74;
end
                default: ;
        endcase*/
			end
	 end
    
endmodule
