//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  10-06-2017                               --
//                                                                       --
//    Fall 2017 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 8                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

// This color mapper is for the background

// color_mapper: Decide which color to be output to VGA for each pixel.
module  color_mapper (input [9:0] DrawX, DrawY, // Current pixel coordinates
                      input [12:0] spriteColor, // for background
							 input [7:0] spriteColor_tracer_1, spriteColor_tracer_2, // for tracer
							 input [7:0] spriteColor_genji_1, spriteColor_genji_2, // for genji
							 input is_tracer_1, is_tracer_2, // current pixel belongs to tracer or not
							 input [23:0] bullet_color_1, bullet_color_2, bullet_color_3, bullet_color_4,
							 input is_healthbar_1, is_healthbar_2, 
							 input [1:0] chara_id_1, chara_id_2,
							 input [9:0] count_k_1, count_k_2, count_l_1, count_l_2, 
							 input is_energybar_1, is_energybar_2,
                      input [23:0] bomb_color_1, bomb_color_2,
							 input [23:0] bullet_show_color_1, bullet_show_color_2,
							 input [7:0] spriteColor_skill,
							 input bomb_warning_color_1, bomb_warning_color_2,
							 input [9:0] bomb_count_1, bomb_count_2,
							 
                      output logic [7:0] VGA_R, VGA_G, VGA_B // VGA RGB output
							 );
    
    logic [7:0] Red, Green, Blue;
    
    // Output colors to VGA
    assign VGA_R = Red;
    assign VGA_G = Green;
    assign VGA_B = Blue;

    // Assign color based on the coordinate
    always_comb
    begin
			if (bullet_show_color_1!=0) begin // not only bullet color
				Red = bullet_show_color_1[23:16];
				Green = bullet_show_color_1[15:8];
				Blue = bullet_show_color_1[7:0];
			end
			else if (bullet_show_color_2!=0) begin
				Red = bullet_show_color_2[23:16];
				Green = bullet_show_color_2[15:8];
				Blue = bullet_show_color_2[7:0];
			end
			else if (is_healthbar_1||is_healthbar_2)
			begin
				Red = 8'h0;
				Green = 8'hff;
				Blue = 8'h0;
			end
			else if (is_energybar_1||is_energybar_2)
			begin
				Red = 8'h0;
				Green = 8'h0;
				Blue = 8'hff;
			end
			else if (bomb_color_1!=24'h0f0f0f) begin
				Red = bomb_color_1[23:16];
				Green = bomb_color_1[15:8];
				Blue = bomb_color_1[7:0];
			end
			else if (bomb_color_2!=24'h0f0f0f) begin
				Red = bomb_color_2[23:16];
				Green = bomb_color_2[15:8];
				Blue = bomb_color_2[7:0];
			end
			else if (bomb_warning_color_1&&bomb_count_1<=10'd19&&bomb_count_1>=10'd0) begin
				Red = 8'hff;
				Green = 8'h99;
				Blue = 8'h33;
			end
			else if (bomb_warning_color_1&&bomb_count_1<=10'd59&&bomb_count_1>=10'd40) begin
				Red = 8'hff;
				Green = 0;
				Blue = 0;
			end
			else if (bomb_warning_color_2&&bomb_count_2<=10'd19&&bomb_count_2>=10'd0) begin
				Red = 8'hff;
				Green = 8'h99;
				Blue = 8'h33;
			end
			else if (bomb_warning_color_2&&bomb_count_2<=10'd59&&bomb_count_2>=10'd40) begin
				Red = 8'hff;
				Green = 0;
				Blue = 0;
			end
			else if (spriteColor_skill!=8'hff) begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_skill)
8'h0:begin Red = 8'h07;Green = 8'h17;Blue = 8'h25;end
8'h1:begin Red = 8'h26;Green = 8'h34;Blue = 8'h40;end
8'h2:begin Red = 8'h27;Green = 8'h35;Blue = 8'h41;end
8'h3:begin Red = 8'h26;Green = 8'h35;Blue = 8'h41;end
8'h4:begin Red = 8'h1a;Green = 8'h29;Blue = 8'h36;end
8'h5:begin Red = 8'h0a;Green = 8'h1a;Blue = 8'h28;end
8'h6:begin Red = 8'h1b;Green = 8'h29;Blue = 8'h36;end
8'h7:begin Red = 8'h1c;Green = 8'h2b;Blue = 8'h38;end
8'h8:begin Red = 8'h22;Green = 8'h30;Blue = 8'h3d;end
8'h9:begin Red = 8'h1f;Green = 8'h2e;Blue = 8'h3a;end
8'ha:begin Red = 8'h09;Green = 8'h19;Blue = 8'h27;end
8'hb:begin Red = 8'h1c;Green = 8'h2a;Blue = 8'h37;end
8'hc:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'hd:begin Red = 8'hfc;Green = 8'hfc;Blue = 8'hfd;end
8'he:begin Red = 8'h21;Green = 8'h30;Blue = 8'h3c;end
8'hf:begin Red = 8'h2e;Green = 8'h3c;Blue = 8'h48;end
8'h10:begin Red = 8'hfe;Green = 8'hfe;Blue = 8'hfe;end
8'h11:begin Red = 8'h1f;Green = 8'h2d;Blue = 8'h3a;end
8'h12:begin Red = 8'hf5;Green = 8'hf6;Blue = 8'hf6;end
8'h13:begin Red = 8'hfa;Green = 8'hfa;Blue = 8'hfa;end
8'h14:begin Red = 8'h22;Green = 8'h31;Blue = 8'h3d;end
8'h15:begin Red = 8'h24;Green = 8'h33;Blue = 8'h3f;end
8'h16:begin Red = 8'h23;Green = 8'h31;Blue = 8'h3e;end
8'h17:begin Red = 8'h1b;Green = 8'h2a;Blue = 8'h37;end
8'h18:begin Red = 8'h1e;Green = 8'h2d;Blue = 8'h3a;end
8'h19:begin Red = 8'h0d;Green = 8'h1c;Blue = 8'h2a;end
8'h1a:begin Red = 8'h25;Green = 8'h33;Blue = 8'h3f;end
8'h1b:begin Red = 8'h26;Green = 8'h34;Blue = 8'h41;end
8'h1c:begin Red = 8'h1e;Green = 8'h2c;Blue = 8'h39;end
8'h1d:begin Red = 8'h25;Green = 8'h33;Blue = 8'h40;end
8'h1e:begin Red = 8'h20;Green = 8'h2e;Blue = 8'h3b;end
8'h1f:begin Red = 8'h1d;Green = 8'h2c;Blue = 8'h39;end
8'h20:begin Red = 8'h0a;Green = 8'h1a;Blue = 8'h27;end
8'h21:begin Red = 8'h25;Green = 8'h32;Blue = 8'h3f;end
8'h22:begin Red = 8'h2a;Green = 8'h37;Blue = 8'h43;end
8'h23:begin Red = 8'h24;Green = 8'h32;Blue = 8'h3f;end
8'h24:begin Red = 8'h20;Green = 8'h2f;Blue = 8'h3b;end
8'h25:begin Red = 8'hf4;Green = 8'hf5;Blue = 8'hf5;end
8'h26:begin Red = 8'hfd;Green = 8'hfd;Blue = 8'hfd;end
8'h27:begin Red = 8'hfa;Green = 8'hfb;Blue = 8'hfb;end
8'h28:begin Red = 8'hfd;Green = 8'hfd;Blue = 8'hfe;end
8'h29:begin Red = 8'hfc;Green = 8'hfc;Blue = 8'hfc;end
8'h2a:begin Red = 8'hf5;Green = 8'hf6;Blue = 8'hf7;end
8'h2b:begin Red = 8'h14;Green = 8'hc9;Blue = 8'hc7;end
8'h2c:begin Red = 8'hef;Green = 8'hf0;Blue = 8'hf1;end
8'h2d:begin Red = 8'hf1;Green = 8'hf2;Blue = 8'hf3;end
8'h2e:begin Red = 8'h1d;Green = 8'h2b;Blue = 8'h38;end
8'h2f:begin Red = 8'h21;Green = 8'h2f;Blue = 8'h3c;end
8'h30:begin Red = 8'h0b;Green = 8'h1b;Blue = 8'h29;end
8'h31:begin Red = 8'h08;Green = 8'h18;Blue = 8'h26;end
8'h32:begin Red = 8'h0e;Green = 8'h1d;Blue = 8'h2b;end
8'h33:begin Red = 8'hf4;Green = 8'hf5;Blue = 8'hf6;end
8'h34:begin Red = 8'h1b;Green = 8'h2a;Blue = 8'h36;end
8'h35:begin Red = 8'h29;Green = 8'h37;Blue = 8'h43;end
8'h36:begin Red = 8'h28;Green = 8'h36;Blue = 8'h42;end
8'h37:begin Red = 8'hf7;Green = 8'hf8;Blue = 8'hf8;end
8'h38:begin Red = 8'h0b;Green = 8'h1a;Blue = 8'h28;end
8'h39:begin Red = 8'h24;Green = 8'h32;Blue = 8'h3e;end
8'h3a:begin Red = 8'hf3;Green = 8'hf4;Blue = 8'hf5;end
8'h3b:begin Red = 8'hf9;Green = 8'hf9;Blue = 8'hf9;end
8'h3c:begin Red = 8'h23;Green = 8'h32;Blue = 8'h3e;end
8'h3d:begin Red = 8'hf9;Green = 8'hf9;Blue = 8'hfa;end
8'h3e:begin Red = 8'h1d;Green = 8'h2c;Blue = 8'h38;end
8'h3f:begin Red = 8'hf0;Green = 8'hf1;Blue = 8'hf2;end
8'h40:begin Red = 8'hf2;Green = 8'hf3;Blue = 8'hf4;end
8'h41:begin Red = 8'h09;Green = 8'h18;Blue = 8'h26;end
8'h42:begin Red = 8'h1c;Green = 8'h2b;Blue = 8'h37;end
8'h43:begin Red = 8'h08;Green = 8'h18;Blue = 8'h25;end
8'h44:begin Red = 8'h0c;Green = 8'h1b;Blue = 8'h29;end
8'h45:begin Red = 8'h19;Green = 8'h28;Blue = 8'h35;end
8'h46:begin Red = 8'h23;Green = 8'h31;Blue = 8'h3d;end
8'h47:begin Red = 8'h16;Green = 8'h30;Blue = 8'h1e;end
8'h48:begin Red = 8'h1b;Green = 8'h35;Blue = 8'h22;end
8'h49:begin Red = 8'h1a;Green = 8'h33;Blue = 8'h21;end
8'h4a:begin Red = 8'h1a;Green = 8'h34;Blue = 8'h22;end
8'h4b:begin Red = 8'h48;Green = 8'h5e;Blue = 8'h49;end
8'h4c:begin Red = 8'h47;Green = 8'h5e;Blue = 8'h49;end
8'h4d:begin Red = 8'h1b;Green = 8'h34;Blue = 8'h22;end
8'h4e:begin Red = 8'h1a;Green = 8'h34;Blue = 8'h21;end
8'h4f:begin Red = 8'h1d;Green = 8'h36;Blue = 8'h24;end
8'h50:begin Red = 8'h17;Green = 8'h30;Blue = 8'h1e;end
8'h51:begin Red = 8'h1d;Green = 8'h36;Blue = 8'h23;end
8'h52:begin Red = 8'h45;Green = 8'h5c;Blue = 8'h47;end
8'h53:begin Red = 8'h1c;Green = 8'h36;Blue = 8'h23;end
8'h54:begin Red = 8'h47;Green = 8'h5d;Blue = 8'h48;end
8'h55:begin Red = 8'h1c;Green = 8'h35;Blue = 8'h23;end
8'h56:begin Red = 8'h45;Green = 8'h5b;Blue = 8'h47;end
8'h57:begin Red = 8'h46;Green = 8'h5d;Blue = 8'h48;end
8'h58:begin Red = 8'h17;Green = 8'h31;Blue = 8'h1f;end
8'h59:begin Red = 8'h18;Green = 8'h31;Blue = 8'h1f;end
8'h5a:begin Red = 8'h46;Green = 8'h5c;Blue = 8'h48;end
8'h5b:begin Red = 8'h2b;Green = 8'h39;Blue = 8'h45;end
8'h5c:begin Red = 8'hf8;Green = 8'hf8;Blue = 8'hf9;end
8'h5d:begin Red = 8'he6;Green = 8'he7;Blue = 8'he9;end
8'h5e:begin Red = 8'h51;Green = 8'h5c;Blue = 8'h66;end
8'h5f:begin Red = 8'hf4;Green = 8'hf4;Blue = 8'hf5;end
8'h60:begin Red = 8'hee;Green = 8'hef;Blue = 8'hf0;end
8'h61:begin Red = 8'hfb;Green = 8'hfb;Blue = 8'hfb;end
8'h62:begin Red = 8'hf7;Green = 8'hf7;Blue = 8'hf8;end
8'h63:begin Red = 8'hdd;Green = 8'hdf;Blue = 8'he1;end
8'h64:begin Red = 8'hd8;Green = 8'hda;Blue = 8'hdd;end
8'h65:begin Red = 8'h3b;Green = 8'h48;Blue = 8'h53;end
8'h66:begin Red = 8'h36;Green = 8'h44;Blue = 8'h4f;end
8'h67:begin Red = 8'h33;Green = 8'h40;Blue = 8'h4c;end
8'h68:begin Red = 8'h2a;Green = 8'h38;Blue = 8'h44;end
8'h69:begin Red = 8'hfd;Green = 8'hfe;Blue = 8'hfe;end
8'h6a:begin Red = 8'hf5;Green = 8'hf5;Blue = 8'hf6;end
8'h6b:begin Red = 8'hed;Green = 8'hee;Blue = 8'hef;end
8'h6c:begin Red = 8'he8;Green = 8'hea;Blue = 8'heb;end
8'h6d:begin Red = 8'h28;Green = 8'h35;Blue = 8'h42;end
8'h6e:begin Red = 8'heb;Green = 8'hec;Blue = 8'hee;end
8'h6f:begin Red = 8'h2c;Green = 8'h3a;Blue = 8'h45;end
8'h70:begin Red = 8'hf8;Green = 8'hf9;Blue = 8'hf9;end
8'h71:begin Red = 8'hf3;Green = 8'hf3;Blue = 8'hf4;end
8'h72:begin Red = 8'he6;Green = 8'he8;Blue = 8'he9;end
8'h73:begin Red = 8'he4;Green = 8'he6;Blue = 8'he8;end
8'h74:begin Red = 8'h0b;Green = 8'h1b;Blue = 8'h28;end
8'h75:begin Red = 8'h46;Green = 8'h5c;Blue = 8'h47;end
8'h76:begin Red = 8'h44;Green = 8'h5b;Blue = 8'h46;end
8'h77:begin Red = 8'h47;Green = 8'h5d;Blue = 8'h49;end
8'h78:begin Red = 8'h44;Green = 8'h5a;Blue = 8'h46;end
8'h79:begin Red = 8'h1d;Green = 8'h37;Blue = 8'h24;end
8'h7a:begin Red = 8'h43;Green = 8'h5a;Blue = 8'h45;end
8'h7b:begin Red = 8'h1e;Green = 8'h37;Blue = 8'h24;end
8'h7c:begin Red = 8'h42;Green = 8'h59;Blue = 8'h45;end
8'h7d:begin Red = 8'h17;Green = 8'h31;Blue = 8'h1e;end
8'h7e:begin Red = 8'h41;Green = 8'h58;Blue = 8'h43;end
8'h7f:begin Red = 8'h40;Green = 8'h57;Blue = 8'h43;end
8'h80:begin Red = 8'h21;Green = 8'h3a;Blue = 8'h27;end
8'h81:begin Red = 8'h20;Green = 8'h39;Blue = 8'h26;end
8'h82:begin Red = 8'h1f;Green = 8'h38;Blue = 8'h26;end
8'h83:begin Red = 8'h1e;Green = 8'h37;Blue = 8'h25;end
8'h84:begin Red = 8'h43;Green = 8'h59;Blue = 8'h45;end
8'h85:begin Red = 8'h25;Green = 8'h3e;Blue = 8'h2b;end
8'h86:begin Red = 8'hfc;Green = 8'hfd;Blue = 8'hfd;end
8'h87:begin Red = 8'hd6;Green = 8'hd9;Blue = 8'hdb;end
8'h88:begin Red = 8'hf6;Green = 8'hf7;Blue = 8'hf7;end
8'h89:begin Red = 8'h2d;Green = 8'h3b;Blue = 8'h47;end
8'h8a:begin Red = 8'h39;Green = 8'h46;Blue = 8'h51;end
8'h8b:begin Red = 8'h0c;Green = 8'h1c;Blue = 8'h29;end
8'h8c:begin Red = 8'hfb;Green = 8'hfb;Blue = 8'hfc;end
8'h8d:begin Red = 8'hfa;Green = 8'hfa;Blue = 8'hfb;end
8'h8e:begin Red = 8'h29;Green = 8'h38;Blue = 8'h44;end
8'h8f:begin Red = 8'h55;Green = 8'h60;Blue = 8'h6a;end
8'h90:begin Red = 8'hcb;Green = 8'hcf;Blue = 8'hd2;end
8'h91:begin Red = 8'he2;Green = 8'he3;Blue = 8'he5;end
8'h92:begin Red = 8'he5;Green = 8'he7;Blue = 8'he8;end
8'h93:begin Red = 8'hf9;Green = 8'hfa;Blue = 8'hfa;end
8'h94:begin Red = 8'hfd;Green = 8'hfc;Blue = 8'hfd;end
8'h95:begin Red = 8'h1f;Green = 8'h2e;Blue = 8'h3b;end
8'h96:begin Red = 8'h25;Green = 8'h34;Blue = 8'h40;end
8'h97:begin Red = 8'h32;Green = 8'h40;Blue = 8'h4b;end
8'h98:begin Red = 8'heb;Green = 8'hed;Blue = 8'hee;end
8'h99:begin Red = 8'hf2;Green = 8'hf3;Blue = 8'hf3;end
8'h9a:begin Red = 8'hbb;Green = 8'hbf;Blue = 8'hc3;end
8'h9b:begin Red = 8'h40;Green = 8'h57;Blue = 8'h42;end
8'h9c:begin Red = 8'h20;Green = 8'h39;Blue = 8'h27;end
8'h9d:begin Red = 8'h26;Green = 8'h3e;Blue = 8'h2c;end
8'h9e:begin Red = 8'h3d;Green = 8'h55;Blue = 8'h40;end
8'h9f:begin Red = 8'h3a;Green = 8'h51;Blue = 8'h3d;end
8'ha0:begin Red = 8'h42;Green = 8'h59;Blue = 8'h44;end
8'ha1:begin Red = 8'h1f;Green = 8'h38;Blue = 8'h25;end
default:;
endcase
			end
			
			
			else if (is_tracer_1&&spriteColor_genji_1!=0)// draw character 1
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_genji_1)
8'h0:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'h1:begin Red = 8'h00;Green = 8'h00;Blue = 8'h00;end
8'h2:begin Red = 8'h15;Green = 8'h15;Blue = 8'h15;end
8'h3:begin Red = 8'h68;Green = 8'h68;Blue = 8'h68;end
8'h4:begin Red = 8'h34;Green = 8'h34;Blue = 8'h34;end
8'h5:begin Red = 8'h38;Green = 8'h38;Blue = 8'h38;end
8'h6:begin Red = 8'h2b;Green = 8'h2b;Blue = 8'h2b;end
8'h7:begin Red = 8'h85;Green = 8'h85;Blue = 8'h85;end
8'h8:begin Red = 8'h89;Green = 8'h89;Blue = 8'h89;end
8'h9:begin Red = 8'h64;Green = 8'h64;Blue = 8'h64;end
8'ha:begin Red = 8'h37;Green = 8'h37;Blue = 8'h37;end
8'hb:begin Red = 8'hd8;Green = 8'hd8;Blue = 8'hd8;end
8'hc:begin Red = 8'h93;Green = 8'hf6;Blue = 8'h5e;end
8'hd:begin Red = 8'h29;Green = 8'h29;Blue = 8'h29;end
8'he:begin Red = 8'hb5;Green = 8'hb5;Blue = 8'hb5;end
8'hf:begin Red = 8'h4b;Green = 8'h4b;Blue = 8'h4b;end
8'h10:begin Red = 8'h3d;Green = 8'h65;Blue = 8'h27;end
8'h11:begin Red = 8'h73;Green = 8'h9d;Blue = 8'h6f;end
8'h12:begin Red = 8'h7a;Green = 8'h5c;Blue = 8'h5c;end
8'h13:begin Red = 8'h34;Green = 8'h36;Blue = 8'h35;end
8'h14:begin Red = 8'h59;Green = 8'h59;Blue = 8'h59;end
8'h15:begin Red = 8'h24;Green = 8'h24;Blue = 8'h24;end
8'h16:begin Red = 8'h89;Green = 8'hfc;Blue = 8'h61;end
8'h17:begin Red = 8'h57;Green = 8'h57;Blue = 8'h57;end
8'h18:begin Red = 8'ha9;Green = 8'hda;Blue = 8'h98;end
8'h19:begin Red = 8'h15;Green = 8'h15;Blue = 8'h17;end
8'h1a:begin Red = 8'h8d;Green = 8'h89;Blue = 8'h88;end
8'h1b:begin Red = 8'h34;Green = 8'h33;Blue = 8'h38;end
8'h1c:begin Red = 8'hda;Green = 8'hdc;Blue = 8'hdb;end
8'h1d:begin Red = 8'h3a;Green = 8'h38;Blue = 8'h38;end
8'h1e:begin Red = 8'h75;Green = 8'h5e;Blue = 8'h66;end
8'h1f:begin Red = 8'hd1;Green = 8'hd1;Blue = 8'hd3;end
8'h20:begin Red = 8'h30;Green = 8'h27;Blue = 8'h2a;end
8'h21:begin Red = 8'h5a;Green = 8'h5b;Blue = 8'h5a;end
8'h22:begin Red = 8'h65;Green = 8'h65;Blue = 8'h67;end
8'h23:begin Red = 8'h7d;Green = 8'h5d;Blue = 8'h5e;end
8'h24:begin Red = 8'h33;Green = 8'h33;Blue = 8'h33;end
8'h25:begin Red = 8'h98;Green = 8'hfd;Blue = 8'h61;end
8'h26:begin Red = 8'h88;Green = 8'h92;Blue = 8'h87;end
8'h27:begin Red = 8'h33;Green = 8'h26;Blue = 8'h27;end
8'h28:begin Red = 8'h35;Green = 8'h64;Blue = 8'h1e;end
8'h29:begin Red = 8'h15;Green = 8'h16;Blue = 8'h16;end
8'h2a:begin Red = 8'h1a;Green = 8'h34;Blue = 8'h36;end
8'h2b:begin Red = 8'hbc;Green = 8'hdf;Blue = 8'h9f;end
8'h2c:begin Red = 8'h32;Green = 8'h32;Blue = 8'h34;end
8'h2d:begin Red = 8'h31;Green = 8'h38;Blue = 8'h31;end
8'h2e:begin Red = 8'h03;Green = 8'h36;Blue = 8'h9b;end
8'h2f:begin Red = 8'hae;Green = 8'hdb;Blue = 8'h96;end
default:;
endcase
			end
			else if (is_tracer_2&&spriteColor_genji_2!=0)// draw character 2
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_genji_2)
8'h0:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'h1:begin Red = 8'h00;Green = 8'h00;Blue = 8'h00;end
8'h2:begin Red = 8'h15;Green = 8'h15;Blue = 8'h15;end
8'h3:begin Red = 8'h68;Green = 8'h68;Blue = 8'h68;end
8'h4:begin Red = 8'h34;Green = 8'h34;Blue = 8'h34;end
8'h5:begin Red = 8'h38;Green = 8'h38;Blue = 8'h38;end
8'h6:begin Red = 8'h2b;Green = 8'h2b;Blue = 8'h2b;end
8'h7:begin Red = 8'h85;Green = 8'h85;Blue = 8'h85;end
8'h8:begin Red = 8'h89;Green = 8'h89;Blue = 8'h89;end
8'h9:begin Red = 8'h64;Green = 8'h64;Blue = 8'h64;end
8'ha:begin Red = 8'h37;Green = 8'h37;Blue = 8'h37;end
8'hb:begin Red = 8'hd8;Green = 8'hd8;Blue = 8'hd8;end
8'hc:begin Red = 8'h93;Green = 8'hf6;Blue = 8'h5e;end
8'hd:begin Red = 8'h29;Green = 8'h29;Blue = 8'h29;end
8'he:begin Red = 8'hb5;Green = 8'hb5;Blue = 8'hb5;end
8'hf:begin Red = 8'h4b;Green = 8'h4b;Blue = 8'h4b;end
8'h10:begin Red = 8'h3d;Green = 8'h65;Blue = 8'h27;end
8'h11:begin Red = 8'h73;Green = 8'h9d;Blue = 8'h6f;end
8'h12:begin Red = 8'h7a;Green = 8'h5c;Blue = 8'h5c;end
8'h13:begin Red = 8'h34;Green = 8'h36;Blue = 8'h35;end
8'h14:begin Red = 8'h59;Green = 8'h59;Blue = 8'h59;end
8'h15:begin Red = 8'h24;Green = 8'h24;Blue = 8'h24;end
8'h16:begin Red = 8'h89;Green = 8'hfc;Blue = 8'h61;end
8'h17:begin Red = 8'h57;Green = 8'h57;Blue = 8'h57;end
8'h18:begin Red = 8'ha9;Green = 8'hda;Blue = 8'h98;end
8'h19:begin Red = 8'h15;Green = 8'h15;Blue = 8'h17;end
8'h1a:begin Red = 8'h8d;Green = 8'h89;Blue = 8'h88;end
8'h1b:begin Red = 8'h34;Green = 8'h33;Blue = 8'h38;end
8'h1c:begin Red = 8'hda;Green = 8'hdc;Blue = 8'hdb;end
8'h1d:begin Red = 8'h3a;Green = 8'h38;Blue = 8'h38;end
8'h1e:begin Red = 8'h75;Green = 8'h5e;Blue = 8'h66;end
8'h1f:begin Red = 8'hd1;Green = 8'hd1;Blue = 8'hd3;end
8'h20:begin Red = 8'h30;Green = 8'h27;Blue = 8'h2a;end
8'h21:begin Red = 8'h5a;Green = 8'h5b;Blue = 8'h5a;end
8'h22:begin Red = 8'h65;Green = 8'h65;Blue = 8'h67;end
8'h23:begin Red = 8'h7d;Green = 8'h5d;Blue = 8'h5e;end
8'h24:begin Red = 8'h33;Green = 8'h33;Blue = 8'h33;end
8'h25:begin Red = 8'h98;Green = 8'hfd;Blue = 8'h61;end
8'h26:begin Red = 8'h88;Green = 8'h92;Blue = 8'h87;end
8'h27:begin Red = 8'h33;Green = 8'h26;Blue = 8'h27;end
8'h28:begin Red = 8'h35;Green = 8'h64;Blue = 8'h1e;end
8'h29:begin Red = 8'h15;Green = 8'h16;Blue = 8'h16;end
8'h2a:begin Red = 8'h1a;Green = 8'h34;Blue = 8'h36;end
8'h2b:begin Red = 8'hbc;Green = 8'hdf;Blue = 8'h9f;end
8'h2c:begin Red = 8'h32;Green = 8'h32;Blue = 8'h34;end
8'h2d:begin Red = 8'h31;Green = 8'h38;Blue = 8'h31;end
8'h2e:begin Red = 8'h03;Green = 8'h36;Blue = 8'h9b;end
8'h2f:begin Red = 8'hae;Green = 8'hdb;Blue = 8'h96;end
default:;
endcase
			end
			else if (is_tracer_1&&spriteColor_tracer_1!=0)// draw character 1
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_tracer_1)
8'h0:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'h1:begin Red = 8'h00;Green = 8'h00;Blue = 8'h00;end
8'h2:begin Red = 8'hfa;Green = 8'hce;Blue = 8'ha8;end
8'h3:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha9;end
8'h4:begin Red = 8'hf2;Green = 8'h9d;Blue = 8'h32;end
8'h5:begin Red = 8'hf1;Green = 8'h9e;Blue = 8'h32;end
8'h6:begin Red = 8'hf3;Green = 8'h7e;Blue = 8'h11;end
8'h7:begin Red = 8'hf3;Green = 8'h9e;Blue = 8'h32;end
8'h8:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha8;end
8'h9:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha8;end
8'ha:begin Red = 8'hf2;Green = 8'h9e;Blue = 8'h33;end
8'hb:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha7;end
8'hc:begin Red = 8'h49;Green = 8'h44;Blue = 8'h40;end
8'hd:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hd0;end
8'he:begin Red = 8'hd7;Green = 8'hd1;Blue = 8'hcf;end
8'hf:begin Red = 8'hd7;Green = 8'hd2;Blue = 8'hd0;end
8'h10:begin Red = 8'hd6;Green = 8'hd0;Blue = 8'hce;end
8'h11:begin Red = 8'h47;Green = 8'h42;Blue = 8'h3f;end
8'h12:begin Red = 8'hfb;Green = 8'hcd;Blue = 8'ha7;end
8'h13:begin Red = 8'h87;Green = 8'h62;Blue = 8'h47;end
8'h14:begin Red = 8'h87;Green = 8'h62;Blue = 8'h46;end
8'h15:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hf1;end
8'h16:begin Red = 8'hd6;Green = 8'hcf;Blue = 8'hcd;end
8'h17:begin Red = 8'hd7;Green = 8'hd0;Blue = 8'hce;end
8'h18:begin Red = 8'h55;Green = 8'h39;Blue = 8'h26;end
8'h19:begin Red = 8'h54;Green = 8'h39;Blue = 8'h25;end
8'h1a:begin Red = 8'h86;Green = 8'h61;Blue = 8'h46;end
8'h1b:begin Red = 8'h87;Green = 8'h62;Blue = 8'h45;end
8'h1c:begin Red = 8'h6a;Green = 8'h66;Blue = 8'h62;end
8'h1d:begin Red = 8'h6c;Green = 8'h66;Blue = 8'h64;end
8'h1e:begin Red = 8'hf1;Green = 8'h9d;Blue = 8'h31;end
8'h1f:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hea;end
8'h20:begin Red = 8'hf3;Green = 8'hee;Blue = 8'heb;end
8'h21:begin Red = 8'hf2;Green = 8'hed;Blue = 8'heb;end
8'h22:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hec;end
8'h23:begin Red = 8'h69;Green = 8'h66;Blue = 8'h61;end
8'h24:begin Red = 8'hbc;Green = 8'hb9;Blue = 8'hbb;end
8'h25:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbd;end
8'h26:begin Red = 8'hbb;Green = 8'hba;Blue = 8'hbc;end
8'h27:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbc;end
8'h28:begin Red = 8'hbc;Green = 8'hb8;Blue = 8'hba;end
8'h29:begin Red = 8'h87;Green = 8'h62;Blue = 8'h48;end
8'h2a:begin Red = 8'h55;Green = 8'h39;Blue = 8'h28;end
8'h2b:begin Red = 8'h54;Green = 8'h39;Blue = 8'h26;end
8'h2c:begin Red = 8'h41;Green = 8'h4f;Blue = 8'h61;end
8'h2d:begin Red = 8'h54;Green = 8'h39;Blue = 8'h28;end
8'h2e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h46;end
8'h2f:begin Red = 8'hf3;Green = 8'hed;Blue = 8'heb;end
8'h30:begin Red = 8'hf4;Green = 8'hed;Blue = 8'heb;end
8'h31:begin Red = 8'hf3;Green = 8'hec;Blue = 8'heb;end
8'h32:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbb;end
8'h33:begin Red = 8'h88;Green = 8'h63;Blue = 8'h47;end
8'h34:begin Red = 8'h55;Green = 8'h39;Blue = 8'h27;end
8'h35:begin Red = 8'h56;Green = 8'h39;Blue = 8'h28;end
8'h36:begin Red = 8'h53;Green = 8'h39;Blue = 8'h25;end
8'h37:begin Red = 8'h55;Green = 8'h38;Blue = 8'h27;end
8'h38:begin Red = 8'h86;Green = 8'h61;Blue = 8'h45;end
8'h39:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd8;end
8'h3a:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd7;end
8'h3b:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd8;end
8'h3c:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd9;end
8'h3d:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd8;end
8'h3e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h48;end
8'h3f:begin Red = 8'h88;Green = 8'h63;Blue = 8'h48;end
8'h40:begin Red = 8'h88;Green = 8'h62;Blue = 8'h47;end
8'h41:begin Red = 8'h6b;Green = 8'h66;Blue = 8'h63;end
8'h42:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd9;end
8'h43:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hd9;end
8'h44:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hda;end
8'h45:begin Red = 8'h86;Green = 8'h61;Blue = 8'h47;end
8'h46:begin Red = 8'h86;Green = 8'h60;Blue = 8'h45;end
8'h47:begin Red = 8'hda;Green = 8'hd8;Blue = 8'hd9;end
8'h48:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd9;end
8'h49:begin Red = 8'h42;Green = 8'h4f;Blue = 8'h61;end
8'h4a:begin Red = 8'h87;Green = 8'h61;Blue = 8'h46;end
8'h4b:begin Red = 8'h87;Green = 8'h61;Blue = 8'h47;end
8'h4c:begin Red = 8'h41;Green = 8'h50;Blue = 8'h62;end
8'h4d:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h44;end
8'h4e:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1c;end
8'h4f:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h22;end
8'h50:begin Red = 8'hf6;Green = 8'h9b;Blue = 8'h11;end
8'h51:begin Red = 8'hf8;Green = 8'h9d;Blue = 8'h14;end
8'h52:begin Red = 8'hf6;Green = 8'h7e;Blue = 8'h18;end
8'h53:begin Red = 8'hf7;Green = 8'h80;Blue = 8'h18;end
8'h54:begin Red = 8'hf3;Green = 8'heb;Blue = 8'he9;end
8'h55:begin Red = 8'hf3;Green = 8'hee;Blue = 8'hec;end
8'h56:begin Red = 8'hf2;Green = 8'heb;Blue = 8'hea;end
8'h57:begin Red = 8'hf3;Green = 8'heb;Blue = 8'hea;end
8'h58:begin Red = 8'hf3;Green = 8'hed;Blue = 8'hea;end
8'h59:begin Red = 8'hd9;Green = 8'hd5;Blue = 8'hd8;end
8'h5a:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1a;end
8'h5b:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h1a;end
8'h5c:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h19;end
8'h5d:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h16;end
8'h5e:begin Red = 8'hfa;Green = 8'hc2;Blue = 8'h1a;end
8'h5f:begin Red = 8'h41;Green = 8'h4e;Blue = 8'h60;end
8'h60:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h17;end
8'h61:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h43;end
8'h62:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h17;end
8'h63:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h43;end
8'h64:begin Red = 8'h42;Green = 8'h51;Blue = 8'h63;end
8'h65:begin Red = 8'hf9;Green = 8'hc2;Blue = 8'h19;end
8'h66:begin Red = 8'hb5;Green = 8'h9a;Blue = 8'h44;end
8'h67:begin Red = 8'h40;Green = 8'h4e;Blue = 8'h60;end
8'h68:begin Red = 8'hb5;Green = 8'h99;Blue = 8'h43;end
8'h69:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h1a;end
8'h6a:begin Red = 8'he2;Green = 8'ha2;Blue = 8'h22;end
8'h6b:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h44;end
8'h6c:begin Red = 8'hf7;Green = 8'h9c;Blue = 8'h14;end
8'h6d:begin Red = 8'hf7;Green = 8'h9b;Blue = 8'h14;end
8'h6e:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h42;end
8'h6f:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h43;end
8'h70:begin Red = 8'hb3;Green = 8'h99;Blue = 8'h43;end
8'h71:begin Red = 8'hf6;Green = 8'h9c;Blue = 8'h14;end
8'h72:begin Red = 8'hf7;Green = 8'h9d;Blue = 8'h14;end
8'h73:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h19;end
8'h74:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h22;end
8'h75:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h20;end
8'h76:begin Red = 8'he0;Green = 8'ha1;Blue = 8'h22;end
8'h77:begin Red = 8'he1;Green = 8'ha3;Blue = 8'h21;end
8'h78:begin Red = 8'hf6;Green = 8'h7d;Blue = 8'h16;end
8'h79:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h23;end
8'h7a:begin Red = 8'hf8;Green = 8'h9e;Blue = 8'h14;end
8'h7b:begin Red = 8'he1;Green = 8'ha1;Blue = 8'h20;end
8'h7c:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h21;end
8'h7d:begin Red = 8'he2;Green = 8'ha4;Blue = 8'h22;end
8'h7e:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h1b;end
8'h7f:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h1a;end
8'h80:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h18;end
8'h81:begin Red = 8'h32;Green = 8'hae;Blue = 8'haf;end
8'h82:begin Red = 8'hfb;Green = 8'hef;Blue = 8'he4;end
8'h83:begin Red = 8'hfc;Green = 8'hef;Blue = 8'he4;end
8'h84:begin Red = 8'hf5;Green = 8'he0;Blue = 8'hbf;end
8'h85:begin Red = 8'hf4;Green = 8'he0;Blue = 8'hbf;end
8'h86:begin Red = 8'hf5;Green = 8'hd6;Blue = 8'hb4;end
8'h87:begin Red = 8'hfb;Green = 8'hef;Blue = 8'he3;end
8'h88:begin Red = 8'h6d;Green = 8'hc4;Blue = 8'hc3;end
8'h89:begin Red = 8'hdd;Green = 8'hd6;Blue = 8'haf;end
8'h8a:begin Red = 8'hdf;Green = 8'hf0;Blue = 8'hf0;end
8'h8b:begin Red = 8'hdf;Green = 8'hf1;Blue = 8'hf0;end
8'h8c:begin Red = 8'hde;Green = 8'hf0;Blue = 8'hf0;end
8'h8d:begin Red = 8'h6b;Green = 8'hc3;Blue = 8'hc3;end
8'h8e:begin Red = 8'hfc;Green = 8'hef;Blue = 8'he3;end
8'h8f:begin Red = 8'h9f;Green = 8'hcd;Blue = 8'hc5;end
8'h90:begin Red = 8'hde;Green = 8'hf0;Blue = 8'hef;end
8'h91:begin Red = 8'h76;Green = 8'hc0;Blue = 8'hbb;end
8'h92:begin Red = 8'h9e;Green = 8'hcd;Blue = 8'hc5;end
8'h93:begin Red = 8'h87;Green = 8'hce;Blue = 8'hce;end
8'h94:begin Red = 8'h89;Green = 8'hce;Blue = 8'hce;end
8'h95:begin Red = 8'hf4;Green = 8'he0;Blue = 8'hbe;end
8'h96:begin Red = 8'hf5;Green = 8'hf9;Blue = 8'hf8;end
8'h97:begin Red = 8'hf5;Green = 8'hfa;Blue = 8'hf9;end
8'h98:begin Red = 8'hf5;Green = 8'hf9;Blue = 8'hf9;end
8'h99:begin Red = 8'h86;Green = 8'hce;Blue = 8'hcd;end
8'h9a:begin Red = 8'hc9;Green = 8'he9;Blue = 8'hea;end
8'h9b:begin Red = 8'hc8;Green = 8'he9;Blue = 8'hea;end
8'h9c:begin Red = 8'hc9;Green = 8'he8;Blue = 8'he9;end
8'h9d:begin Red = 8'h9f;Green = 8'hcd;Blue = 8'hc6;end
8'h9e:begin Red = 8'h76;Green = 8'hc0;Blue = 8'hbc;end
8'h9f:begin Red = 8'h66;Green = 8'hc7;Blue = 8'hcd;end
8'ha0:begin Red = 8'hf6;Green = 8'hf9;Blue = 8'hf9;end
8'ha1:begin Red = 8'h77;Green = 8'hc0;Blue = 8'hbc;end
8'ha2:begin Red = 8'h75;Green = 8'hc0;Blue = 8'hbb;end
8'ha3:begin Red = 8'he0;Green = 8'hf2;Blue = 8'hf3;end
8'ha4:begin Red = 8'he0;Green = 8'hf2;Blue = 8'hf2;end
8'ha5:begin Red = 8'he1;Green = 8'hf2;Blue = 8'hf3;end
8'ha6:begin Red = 8'h88;Green = 8'hce;Blue = 8'hce;end
8'ha7:begin Red = 8'he0;Green = 8'hf3;Blue = 8'hf3;end
8'ha8:begin Red = 8'h9e;Green = 8'hcc;Blue = 8'hc5;end
8'ha9:begin Red = 8'he1;Green = 8'hf3;Blue = 8'hf3;end
8'haa:begin Red = 8'h67;Green = 8'hc7;Blue = 8'hcd;end
8'hab:begin Red = 8'h66;Green = 8'hc7;Blue = 8'hce;end
8'hac:begin Red = 8'hc3;Green = 8'hdf;Blue = 8'hc4;end
8'had:begin Red = 8'hfa;Green = 8'heb;Blue = 8'hb8;end
8'hae:begin Red = 8'he7;Green = 8'he1;Blue = 8'hba;end
8'haf:begin Red = 8'hf8;Green = 8'hdf;Blue = 8'hb4;end
8'hb0:begin Red = 8'hf9;Green = 8'he0;Blue = 8'hb5;end
8'hb1:begin Red = 8'hf8;Green = 8'hd6;Blue = 8'hb7;end
8'hb2:begin Red = 8'hf9;Green = 8'hd7;Blue = 8'hb7;end
8'hb3:begin Red = 8'hfa;Green = 8'heb;Blue = 8'hb7;end
8'hb4:begin Red = 8'hfb;Green = 8'heb;Blue = 8'hb7;end
8'hb5:begin Red = 8'hfa;Green = 8'heb;Blue = 8'hb6;end
8'hb6:begin Red = 8'hfb;Green = 8'hec;Blue = 8'hb7;end
8'hb7:begin Red = 8'hc2;Green = 8'hde;Blue = 8'hc4;end
8'hb8:begin Red = 8'hfb;Green = 8'heb;Blue = 8'hb6;end
8'hb9:begin Red = 8'h67;Green = 8'hc8;Blue = 8'hce;end
8'hba:begin Red = 8'hfa;Green = 8'hec;Blue = 8'hb7;end
8'hbb:begin Red = 8'hc4;Green = 8'hdf;Blue = 8'hc4;end
8'hbc:begin Red = 8'h65;Green = 8'hc7;Blue = 8'hcd;end
8'hbd:begin Red = 8'he8;Green = 8'he1;Blue = 8'hba;end
8'hbe:begin Red = 8'hf9;Green = 8'hdf;Blue = 8'hb5;end
8'hbf:begin Red = 8'hc2;Green = 8'hdf;Blue = 8'hc4;end
8'hc0:begin Red = 8'hf8;Green = 8'he0;Blue = 8'hb5;end
8'hc1:begin Red = 8'hf9;Green = 8'hd6;Blue = 8'hb7;end
8'hc2:begin Red = 8'he8;Green = 8'he2;Blue = 8'hba;end
8'hc3:begin Red = 8'he7;Green = 8'he1;Blue = 8'hb9;end
8'hc4:begin Red = 8'he6;Green = 8'he1;Blue = 8'hba;end
8'hc5:begin Red = 8'he7;Green = 8'he2;Blue = 8'hb9;end
8'hc6:begin Red = 8'hf8;Green = 8'hd6;Blue = 8'hb6;end
8'hc7:begin Red = 8'hb4;Green = 8'h77;Blue = 8'hff;end
8'hc8:begin Red = 8'hfe;Green = 8'he5;Blue = 8'hff;end
8'hc9:begin Red = 8'hfb;Green = 8'hcb;Blue = 8'hff;end
8'hca:begin Red = 8'hfb;Green = 8'hba;Blue = 8'hff;end
8'hcb:begin Red = 8'hfe;Green = 8'he4;Blue = 8'hff;end
8'hcc:begin Red = 8'hc9;Green = 8'h9b;Blue = 8'hff;end
8'hcd:begin Red = 8'hf3;Green = 8'hba;Blue = 8'hff;end
8'hce:begin Red = 8'hf3;Green = 8'he6;Blue = 8'hff;end
8'hcf:begin Red = 8'hf3;Green = 8'he7;Blue = 8'hff;end
8'hd0:begin Red = 8'hc9;Green = 8'h9a;Blue = 8'hff;end
8'hd1:begin Red = 8'hdc;Green = 8'hab;Blue = 8'hff;end
8'hd2:begin Red = 8'hf3;Green = 8'hbb;Blue = 8'hff;end
8'hd3:begin Red = 8'hf3;Green = 8'he5;Blue = 8'hff;end
8'hd4:begin Red = 8'hcd;Green = 8'h95;Blue = 8'hff;end
8'hd5:begin Red = 8'hdb;Green = 8'hab;Blue = 8'hff;end
8'hd6:begin Red = 8'hd3;Green = 8'had;Blue = 8'hff;end
8'hd7:begin Red = 8'hd4;Green = 8'had;Blue = 8'hff;end
8'hd8:begin Red = 8'hfb;Green = 8'hf5;Blue = 8'hff;end
8'hd9:begin Red = 8'hfb;Green = 8'hf6;Blue = 8'hff;end
8'hda:begin Red = 8'heb;Green = 8'hda;Blue = 8'hff;end
8'hdb:begin Red = 8'heb;Green = 8'hd9;Blue = 8'hff;end
8'hdc:begin Red = 8'hc7;Green = 8'ha1;Blue = 8'hff;end
8'hdd:begin Red = 8'hdc;Green = 8'hac;Blue = 8'hff;end
8'hde:begin Red = 8'hfc;Green = 8'hf5;Blue = 8'hff;end
8'hdf:begin Red = 8'hcc;Green = 8'h95;Blue = 8'hff;end
8'he0:begin Red = 8'hf4;Green = 8'hea;Blue = 8'hff;end
8'he1:begin Red = 8'hf4;Green = 8'he9;Blue = 8'hff;end
8'he2:begin Red = 8'hdb;Green = 8'haa;Blue = 8'hff;end
8'he3:begin Red = 8'hc7;Green = 8'ha2;Blue = 8'hff;end
8'he4:begin Red = 8'he9;Green = 8'hc9;Blue = 8'hff;end
8'he5:begin Red = 8'hfd;Green = 8'hde;Blue = 8'hff;end
8'he6:begin Red = 8'hf6;Green = 8'hcd;Blue = 8'hff;end
8'he7:begin Red = 8'hfc;Green = 8'hca;Blue = 8'hff;end
8'he8:begin Red = 8'hfd;Green = 8'hcb;Blue = 8'hff;end
8'he9:begin Red = 8'hfc;Green = 8'hba;Blue = 8'hff;end
8'hea:begin Red = 8'hfd;Green = 8'hbb;Blue = 8'hff;end
8'heb:begin Red = 8'hfb;Green = 8'hf4;Blue = 8'hff;end
8'hec:begin Red = 8'hfe;Green = 8'hde;Blue = 8'hff;end
8'hed:begin Red = 8'hfd;Green = 8'hdd;Blue = 8'hff;end
8'hee:begin Red = 8'he9;Green = 8'hc8;Blue = 8'hff;end
8'hef:begin Red = 8'hfd;Green = 8'hca;Blue = 8'hff;end
8'hf0:begin Red = 8'hf6;Green = 8'hce;Blue = 8'hff;end
8'hf1:begin Red = 8'hfc;Green = 8'hbb;Blue = 8'hff;end

endcase
			end
			else if (is_tracer_2&&spriteColor_tracer_2!=0) // draw character 2
			begin
				Red = 8'hff;
				Green = 8'hff;
				Blue = 8'hff;
case(spriteColor_tracer_2)
8'h0:begin Red = 8'hff;Green = 8'hff;Blue = 8'hff;end
8'h1:begin Red = 8'h00;Green = 8'h00;Blue = 8'h00;end
8'h2:begin Red = 8'hfa;Green = 8'hce;Blue = 8'ha8;end
8'h3:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha9;end
8'h4:begin Red = 8'hf2;Green = 8'h9d;Blue = 8'h32;end
8'h5:begin Red = 8'hf1;Green = 8'h9e;Blue = 8'h32;end
8'h6:begin Red = 8'hf3;Green = 8'h7e;Blue = 8'h11;end
8'h7:begin Red = 8'hf3;Green = 8'h9e;Blue = 8'h32;end
8'h8:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha8;end
8'h9:begin Red = 8'hfb;Green = 8'hce;Blue = 8'ha8;end
8'ha:begin Red = 8'hf2;Green = 8'h9e;Blue = 8'h33;end
8'hb:begin Red = 8'hfa;Green = 8'hcd;Blue = 8'ha7;end
8'hc:begin Red = 8'h49;Green = 8'h44;Blue = 8'h40;end
8'hd:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hd0;end
8'he:begin Red = 8'hd7;Green = 8'hd1;Blue = 8'hcf;end
8'hf:begin Red = 8'hd7;Green = 8'hd2;Blue = 8'hd0;end
8'h10:begin Red = 8'hd6;Green = 8'hd0;Blue = 8'hce;end
8'h11:begin Red = 8'h47;Green = 8'h42;Blue = 8'h3f;end
8'h12:begin Red = 8'hfb;Green = 8'hcd;Blue = 8'ha7;end
8'h13:begin Red = 8'h87;Green = 8'h62;Blue = 8'h47;end
8'h14:begin Red = 8'h87;Green = 8'h62;Blue = 8'h46;end
8'h15:begin Red = 8'h0d;Green = 8'h57;Blue = 8'hf1;end
8'h16:begin Red = 8'hd6;Green = 8'hcf;Blue = 8'hcd;end
8'h17:begin Red = 8'hd7;Green = 8'hd0;Blue = 8'hce;end
8'h18:begin Red = 8'h55;Green = 8'h39;Blue = 8'h26;end
8'h19:begin Red = 8'h54;Green = 8'h39;Blue = 8'h25;end
8'h1a:begin Red = 8'h86;Green = 8'h61;Blue = 8'h46;end
8'h1b:begin Red = 8'h87;Green = 8'h62;Blue = 8'h45;end
8'h1c:begin Red = 8'h6a;Green = 8'h66;Blue = 8'h62;end
8'h1d:begin Red = 8'h6c;Green = 8'h66;Blue = 8'h64;end
8'h1e:begin Red = 8'hf1;Green = 8'h9d;Blue = 8'h31;end
8'h1f:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hea;end
8'h20:begin Red = 8'hf3;Green = 8'hee;Blue = 8'heb;end
8'h21:begin Red = 8'hf2;Green = 8'hed;Blue = 8'heb;end
8'h22:begin Red = 8'hf3;Green = 8'hec;Blue = 8'hec;end
8'h23:begin Red = 8'h69;Green = 8'h66;Blue = 8'h61;end
8'h24:begin Red = 8'hbc;Green = 8'hb9;Blue = 8'hbb;end
8'h25:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbd;end
8'h26:begin Red = 8'hbb;Green = 8'hba;Blue = 8'hbc;end
8'h27:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbc;end
8'h28:begin Red = 8'hbc;Green = 8'hb8;Blue = 8'hba;end
8'h29:begin Red = 8'h87;Green = 8'h62;Blue = 8'h48;end
8'h2a:begin Red = 8'h55;Green = 8'h39;Blue = 8'h28;end
8'h2b:begin Red = 8'h54;Green = 8'h39;Blue = 8'h26;end
8'h2c:begin Red = 8'h41;Green = 8'h4f;Blue = 8'h61;end
8'h2d:begin Red = 8'h54;Green = 8'h39;Blue = 8'h28;end
8'h2e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h46;end
8'h2f:begin Red = 8'hf3;Green = 8'hed;Blue = 8'heb;end
8'h30:begin Red = 8'hf4;Green = 8'hed;Blue = 8'heb;end
8'h31:begin Red = 8'hf3;Green = 8'hec;Blue = 8'heb;end
8'h32:begin Red = 8'hbc;Green = 8'hba;Blue = 8'hbb;end
8'h33:begin Red = 8'h88;Green = 8'h63;Blue = 8'h47;end
8'h34:begin Red = 8'h55;Green = 8'h39;Blue = 8'h27;end
8'h35:begin Red = 8'h56;Green = 8'h39;Blue = 8'h28;end
8'h36:begin Red = 8'h53;Green = 8'h39;Blue = 8'h25;end
8'h37:begin Red = 8'h55;Green = 8'h38;Blue = 8'h27;end
8'h38:begin Red = 8'h86;Green = 8'h61;Blue = 8'h45;end
8'h39:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd8;end
8'h3a:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd7;end
8'h3b:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd8;end
8'h3c:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd9;end
8'h3d:begin Red = 8'hd9;Green = 8'hd6;Blue = 8'hd8;end
8'h3e:begin Red = 8'h87;Green = 8'h63;Blue = 8'h48;end
8'h3f:begin Red = 8'h88;Green = 8'h63;Blue = 8'h48;end
8'h40:begin Red = 8'h88;Green = 8'h62;Blue = 8'h47;end
8'h41:begin Red = 8'h6b;Green = 8'h66;Blue = 8'h63;end
8'h42:begin Red = 8'hda;Green = 8'hd7;Blue = 8'hd9;end
8'h43:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hd9;end
8'h44:begin Red = 8'hd9;Green = 8'hd8;Blue = 8'hda;end
8'h45:begin Red = 8'h86;Green = 8'h61;Blue = 8'h47;end
8'h46:begin Red = 8'h86;Green = 8'h60;Blue = 8'h45;end
8'h47:begin Red = 8'hda;Green = 8'hd8;Blue = 8'hd9;end
8'h48:begin Red = 8'hd9;Green = 8'hd7;Blue = 8'hd9;end
8'h49:begin Red = 8'h42;Green = 8'h4f;Blue = 8'h61;end
8'h4a:begin Red = 8'h87;Green = 8'h61;Blue = 8'h46;end
8'h4b:begin Red = 8'h87;Green = 8'h61;Blue = 8'h47;end
8'h4c:begin Red = 8'h41;Green = 8'h50;Blue = 8'h62;end
8'h4d:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h44;end
8'h4e:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1c;end
8'h4f:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h22;end
8'h50:begin Red = 8'hf6;Green = 8'h9b;Blue = 8'h11;end
8'h51:begin Red = 8'hf8;Green = 8'h9d;Blue = 8'h14;end
8'h52:begin Red = 8'hf6;Green = 8'h7e;Blue = 8'h18;end
8'h53:begin Red = 8'hf7;Green = 8'h80;Blue = 8'h18;end
8'h54:begin Red = 8'hf3;Green = 8'heb;Blue = 8'he9;end
8'h55:begin Red = 8'hf3;Green = 8'hee;Blue = 8'hec;end
8'h56:begin Red = 8'hf2;Green = 8'heb;Blue = 8'hea;end
8'h57:begin Red = 8'hf3;Green = 8'heb;Blue = 8'hea;end
8'h58:begin Red = 8'hf3;Green = 8'hed;Blue = 8'hea;end
8'h59:begin Red = 8'hd9;Green = 8'hd5;Blue = 8'hd8;end
8'h5a:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h1a;end
8'h5b:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h1a;end
8'h5c:begin Red = 8'hf9;Green = 8'hc1;Blue = 8'h19;end
8'h5d:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h16;end
8'h5e:begin Red = 8'hfa;Green = 8'hc2;Blue = 8'h1a;end
8'h5f:begin Red = 8'h41;Green = 8'h4e;Blue = 8'h60;end
8'h60:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h17;end
8'h61:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h43;end
8'h62:begin Red = 8'hfa;Green = 8'hc1;Blue = 8'h17;end
8'h63:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h43;end
8'h64:begin Red = 8'h42;Green = 8'h51;Blue = 8'h63;end
8'h65:begin Red = 8'hf9;Green = 8'hc2;Blue = 8'h19;end
8'h66:begin Red = 8'hb5;Green = 8'h9a;Blue = 8'h44;end
8'h67:begin Red = 8'h40;Green = 8'h4e;Blue = 8'h60;end
8'h68:begin Red = 8'hb5;Green = 8'h99;Blue = 8'h43;end
8'h69:begin Red = 8'hf9;Green = 8'hc0;Blue = 8'h1a;end
8'h6a:begin Red = 8'he2;Green = 8'ha2;Blue = 8'h22;end
8'h6b:begin Red = 8'hb4;Green = 8'h99;Blue = 8'h44;end
8'h6c:begin Red = 8'hf7;Green = 8'h9c;Blue = 8'h14;end
8'h6d:begin Red = 8'hf7;Green = 8'h9b;Blue = 8'h14;end
8'h6e:begin Red = 8'hb3;Green = 8'h98;Blue = 8'h42;end
8'h6f:begin Red = 8'hb4;Green = 8'h9a;Blue = 8'h43;end
8'h70:begin Red = 8'hb3;Green = 8'h99;Blue = 8'h43;end
8'h71:begin Red = 8'hf6;Green = 8'h9c;Blue = 8'h14;end
8'h72:begin Red = 8'hf7;Green = 8'h9d;Blue = 8'h14;end
8'h73:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h19;end
8'h74:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h22;end
8'h75:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h20;end
8'h76:begin Red = 8'he0;Green = 8'ha1;Blue = 8'h22;end
8'h77:begin Red = 8'he1;Green = 8'ha3;Blue = 8'h21;end
8'h78:begin Red = 8'hf6;Green = 8'h7d;Blue = 8'h16;end
8'h79:begin Red = 8'he2;Green = 8'ha3;Blue = 8'h23;end
8'h7a:begin Red = 8'hf8;Green = 8'h9e;Blue = 8'h14;end
8'h7b:begin Red = 8'he1;Green = 8'ha1;Blue = 8'h20;end
8'h7c:begin Red = 8'he1;Green = 8'ha2;Blue = 8'h21;end
8'h7d:begin Red = 8'he2;Green = 8'ha4;Blue = 8'h22;end
8'h7e:begin Red = 8'hf7;Green = 8'h7f;Blue = 8'h1b;end
8'h7f:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h1a;end
8'h80:begin Red = 8'hf6;Green = 8'h7f;Blue = 8'h18;end
8'h81:begin Red = 8'h32;Green = 8'hae;Blue = 8'haf;end
8'h82:begin Red = 8'hfb;Green = 8'hef;Blue = 8'he4;end
8'h83:begin Red = 8'hfc;Green = 8'hef;Blue = 8'he4;end
8'h84:begin Red = 8'hf5;Green = 8'he0;Blue = 8'hbf;end
8'h85:begin Red = 8'hf4;Green = 8'he0;Blue = 8'hbf;end
8'h86:begin Red = 8'hf5;Green = 8'hd6;Blue = 8'hb4;end
8'h87:begin Red = 8'hfb;Green = 8'hef;Blue = 8'he3;end
8'h88:begin Red = 8'h6d;Green = 8'hc4;Blue = 8'hc3;end
8'h89:begin Red = 8'hdd;Green = 8'hd6;Blue = 8'haf;end
8'h8a:begin Red = 8'hdf;Green = 8'hf0;Blue = 8'hf0;end
8'h8b:begin Red = 8'hdf;Green = 8'hf1;Blue = 8'hf0;end
8'h8c:begin Red = 8'hde;Green = 8'hf0;Blue = 8'hf0;end
8'h8d:begin Red = 8'h6b;Green = 8'hc3;Blue = 8'hc3;end
8'h8e:begin Red = 8'hfc;Green = 8'hef;Blue = 8'he3;end
8'h8f:begin Red = 8'h9f;Green = 8'hcd;Blue = 8'hc5;end
8'h90:begin Red = 8'hde;Green = 8'hf0;Blue = 8'hef;end
8'h91:begin Red = 8'h76;Green = 8'hc0;Blue = 8'hbb;end
8'h92:begin Red = 8'h9e;Green = 8'hcd;Blue = 8'hc5;end
8'h93:begin Red = 8'h87;Green = 8'hce;Blue = 8'hce;end
8'h94:begin Red = 8'h89;Green = 8'hce;Blue = 8'hce;end
8'h95:begin Red = 8'hf4;Green = 8'he0;Blue = 8'hbe;end
8'h96:begin Red = 8'hf5;Green = 8'hf9;Blue = 8'hf8;end
8'h97:begin Red = 8'hf5;Green = 8'hfa;Blue = 8'hf9;end
8'h98:begin Red = 8'hf5;Green = 8'hf9;Blue = 8'hf9;end
8'h99:begin Red = 8'h86;Green = 8'hce;Blue = 8'hcd;end
8'h9a:begin Red = 8'hc9;Green = 8'he9;Blue = 8'hea;end
8'h9b:begin Red = 8'hc8;Green = 8'he9;Blue = 8'hea;end
8'h9c:begin Red = 8'hc9;Green = 8'he8;Blue = 8'he9;end
8'h9d:begin Red = 8'h9f;Green = 8'hcd;Blue = 8'hc6;end
8'h9e:begin Red = 8'h76;Green = 8'hc0;Blue = 8'hbc;end
8'h9f:begin Red = 8'h66;Green = 8'hc7;Blue = 8'hcd;end
8'ha0:begin Red = 8'hf6;Green = 8'hf9;Blue = 8'hf9;end
8'ha1:begin Red = 8'h77;Green = 8'hc0;Blue = 8'hbc;end
8'ha2:begin Red = 8'h75;Green = 8'hc0;Blue = 8'hbb;end
8'ha3:begin Red = 8'he0;Green = 8'hf2;Blue = 8'hf3;end
8'ha4:begin Red = 8'he0;Green = 8'hf2;Blue = 8'hf2;end
8'ha5:begin Red = 8'he1;Green = 8'hf2;Blue = 8'hf3;end
8'ha6:begin Red = 8'h88;Green = 8'hce;Blue = 8'hce;end
8'ha7:begin Red = 8'he0;Green = 8'hf3;Blue = 8'hf3;end
8'ha8:begin Red = 8'h9e;Green = 8'hcc;Blue = 8'hc5;end
8'ha9:begin Red = 8'he1;Green = 8'hf3;Blue = 8'hf3;end
8'haa:begin Red = 8'h67;Green = 8'hc7;Blue = 8'hcd;end
8'hab:begin Red = 8'h66;Green = 8'hc7;Blue = 8'hce;end
8'hac:begin Red = 8'hc3;Green = 8'hdf;Blue = 8'hc4;end
8'had:begin Red = 8'hfa;Green = 8'heb;Blue = 8'hb8;end
8'hae:begin Red = 8'he7;Green = 8'he1;Blue = 8'hba;end
8'haf:begin Red = 8'hf8;Green = 8'hdf;Blue = 8'hb4;end
8'hb0:begin Red = 8'hf9;Green = 8'he0;Blue = 8'hb5;end
8'hb1:begin Red = 8'hf8;Green = 8'hd6;Blue = 8'hb7;end
8'hb2:begin Red = 8'hf9;Green = 8'hd7;Blue = 8'hb7;end
8'hb3:begin Red = 8'hfa;Green = 8'heb;Blue = 8'hb7;end
8'hb4:begin Red = 8'hfb;Green = 8'heb;Blue = 8'hb7;end
8'hb5:begin Red = 8'hfa;Green = 8'heb;Blue = 8'hb6;end
8'hb6:begin Red = 8'hfb;Green = 8'hec;Blue = 8'hb7;end
8'hb7:begin Red = 8'hc2;Green = 8'hde;Blue = 8'hc4;end
8'hb8:begin Red = 8'hfb;Green = 8'heb;Blue = 8'hb6;end
8'hb9:begin Red = 8'h67;Green = 8'hc8;Blue = 8'hce;end
8'hba:begin Red = 8'hfa;Green = 8'hec;Blue = 8'hb7;end
8'hbb:begin Red = 8'hc4;Green = 8'hdf;Blue = 8'hc4;end
8'hbc:begin Red = 8'h65;Green = 8'hc7;Blue = 8'hcd;end
8'hbd:begin Red = 8'he8;Green = 8'he1;Blue = 8'hba;end
8'hbe:begin Red = 8'hf9;Green = 8'hdf;Blue = 8'hb5;end
8'hbf:begin Red = 8'hc2;Green = 8'hdf;Blue = 8'hc4;end
8'hc0:begin Red = 8'hf8;Green = 8'he0;Blue = 8'hb5;end
8'hc1:begin Red = 8'hf9;Green = 8'hd6;Blue = 8'hb7;end
8'hc2:begin Red = 8'he8;Green = 8'he2;Blue = 8'hba;end
8'hc3:begin Red = 8'he7;Green = 8'he1;Blue = 8'hb9;end
8'hc4:begin Red = 8'he6;Green = 8'he1;Blue = 8'hba;end
8'hc5:begin Red = 8'he7;Green = 8'he2;Blue = 8'hb9;end
8'hc6:begin Red = 8'hf8;Green = 8'hd6;Blue = 8'hb6;end
8'hc7:begin Red = 8'hb4;Green = 8'h77;Blue = 8'hff;end
8'hc8:begin Red = 8'hfe;Green = 8'he5;Blue = 8'hff;end
8'hc9:begin Red = 8'hfb;Green = 8'hcb;Blue = 8'hff;end
8'hca:begin Red = 8'hfb;Green = 8'hba;Blue = 8'hff;end
8'hcb:begin Red = 8'hfe;Green = 8'he4;Blue = 8'hff;end
8'hcc:begin Red = 8'hc9;Green = 8'h9b;Blue = 8'hff;end
8'hcd:begin Red = 8'hf3;Green = 8'hba;Blue = 8'hff;end
8'hce:begin Red = 8'hf3;Green = 8'he6;Blue = 8'hff;end
8'hcf:begin Red = 8'hf3;Green = 8'he7;Blue = 8'hff;end
8'hd0:begin Red = 8'hc9;Green = 8'h9a;Blue = 8'hff;end
8'hd1:begin Red = 8'hdc;Green = 8'hab;Blue = 8'hff;end
8'hd2:begin Red = 8'hf3;Green = 8'hbb;Blue = 8'hff;end
8'hd3:begin Red = 8'hf3;Green = 8'he5;Blue = 8'hff;end
8'hd4:begin Red = 8'hcd;Green = 8'h95;Blue = 8'hff;end
8'hd5:begin Red = 8'hdb;Green = 8'hab;Blue = 8'hff;end
8'hd6:begin Red = 8'hd3;Green = 8'had;Blue = 8'hff;end
8'hd7:begin Red = 8'hd4;Green = 8'had;Blue = 8'hff;end
8'hd8:begin Red = 8'hfb;Green = 8'hf5;Blue = 8'hff;end
8'hd9:begin Red = 8'hfb;Green = 8'hf6;Blue = 8'hff;end
8'hda:begin Red = 8'heb;Green = 8'hda;Blue = 8'hff;end
8'hdb:begin Red = 8'heb;Green = 8'hd9;Blue = 8'hff;end
8'hdc:begin Red = 8'hc7;Green = 8'ha1;Blue = 8'hff;end
8'hdd:begin Red = 8'hdc;Green = 8'hac;Blue = 8'hff;end
8'hde:begin Red = 8'hfc;Green = 8'hf5;Blue = 8'hff;end
8'hdf:begin Red = 8'hcc;Green = 8'h95;Blue = 8'hff;end
8'he0:begin Red = 8'hf4;Green = 8'hea;Blue = 8'hff;end
8'he1:begin Red = 8'hf4;Green = 8'he9;Blue = 8'hff;end
8'he2:begin Red = 8'hdb;Green = 8'haa;Blue = 8'hff;end
8'he3:begin Red = 8'hc7;Green = 8'ha2;Blue = 8'hff;end
8'he4:begin Red = 8'he9;Green = 8'hc9;Blue = 8'hff;end
8'he5:begin Red = 8'hfd;Green = 8'hde;Blue = 8'hff;end
8'he6:begin Red = 8'hf6;Green = 8'hcd;Blue = 8'hff;end
8'he7:begin Red = 8'hfc;Green = 8'hca;Blue = 8'hff;end
8'he8:begin Red = 8'hfd;Green = 8'hcb;Blue = 8'hff;end
8'he9:begin Red = 8'hfc;Green = 8'hba;Blue = 8'hff;end
8'hea:begin Red = 8'hfd;Green = 8'hbb;Blue = 8'hff;end
8'heb:begin Red = 8'hfb;Green = 8'hf4;Blue = 8'hff;end
8'hec:begin Red = 8'hfe;Green = 8'hde;Blue = 8'hff;end
8'hed:begin Red = 8'hfd;Green = 8'hdd;Blue = 8'hff;end
8'hee:begin Red = 8'he9;Green = 8'hc8;Blue = 8'hff;end
8'hef:begin Red = 8'hfd;Green = 8'hca;Blue = 8'hff;end
8'hf0:begin Red = 8'hf6;Green = 8'hce;Blue = 8'hff;end
8'hf1:begin Red = 8'hfc;Green = 8'hbb;Blue = 8'hff;end

endcase
			end
			else if (bullet_color_3!=24'h000000) begin
					Red = bullet_color_3[23:16];
					Green = bullet_color_3[15:8];
					Blue = bullet_color_3[7:0];
			end
			else if (bullet_color_4!=24'h000000) begin
					Red = bullet_color_4[23:16];
					Green = bullet_color_4[15:8];
					Blue = bullet_color_4[7:0];
			end
			else if (bullet_color_1!=24'h000000) begin // draw bullet
					Red = bullet_color_1[23:16];
					Green = bullet_color_1[15:8];
					Blue = bullet_color_1[7:0];
			end
			else if (bullet_color_2!=24'h000000) begin
					Red = bullet_color_2[23:16];
					Green = bullet_color_2[15:8];
					Blue = bullet_color_2[7:0];
			end
			else // draw background
			begin
				  Red   = 8'h80;
				  Green = 8'h80;
				  Blue  = 8'h80;/*
				  case(spriteColor)
13'h0:    begin Red = 8'h64;    Green = 8'h7b;    Blue = 8'h81;
end 13'h1:    begin Red = 8'h66;    Green = 8'h7d;    Blue = 8'h84;
end 13'h2:    begin Red = 8'h55;    Green = 8'h6a;    Blue = 8'h70;
end 13'h3:    begin Red = 8'h5a;    Green = 8'h6f;    Blue = 8'h75;
end 13'h4:    begin Red = 8'h56;    Green = 8'h6e;    Blue = 8'h77;
end 13'h5:    begin Red = 8'ha1;    Green = 8'hf7;    Blue = 8'hff;
end 13'h6:    begin Red = 8'h9b;    Green = 8'he3;    Blue = 8'hf9;
end 13'h7:    begin Red = 8'h90;    Green = 8'he2;    Blue = 8'hea;
end 13'h8:    begin Red = 8'h8e;    Green = 8'hcd;    Blue = 8'he5;
end 13'h9:    begin Red = 8'h90;    Green = 8'hce;    Blue = 8'hdf;
end 13'ha:    begin Red = 8'h91;    Green = 8'hda;    Blue = 8'hed;
end 13'hb:    begin Red = 8'h95;    Green = 8'hd9;    Blue = 8'hed;
end 13'hc:    begin Red = 8'h94;    Green = 8'he2;    Blue = 8'hfb;
end 13'hd:    begin Red = 8'h80;    Green = 8'h98;    Blue = 8'h94;
end 13'he:    begin Red = 8'h84;    Green = 8'h9b;    Blue = 8'ha0;
end 13'hf:    begin Red = 8'h75;    Green = 8'h9a;    Blue = 8'h92;
end 13'h10:    begin Red = 8'h7f;    Green = 8'h97;    Blue = 8'h98;
end 13'h11:    begin Red = 8'h7d;    Green = 8'h95;    Blue = 8'h97;
end 13'h12:    begin Red = 8'h82;    Green = 8'h9a;    Blue = 8'h9b;
end 13'h13:    begin Red = 8'h5c;    Green = 8'h73;    Blue = 8'h79;
end 13'h14:    begin Red = 8'h61;    Green = 8'h78;    Blue = 8'h7f;
end 13'h15:    begin Red = 8'h65;    Green = 8'h7e;    Blue = 8'h87;
end 13'h16:    begin Red = 8'h52;    Green = 8'h60;    Blue = 8'h66;
end 13'h17:    begin Red = 8'h58;    Green = 8'h67;    Blue = 8'h6c;
end 13'h18:    begin Red = 8'h55;    Green = 8'h65;    Blue = 8'h69;
end 13'h19:    begin Red = 8'h54;    Green = 8'h55;    Blue = 8'h61;
end 13'h1a:    begin Red = 8'h8e;    Green = 8'hcf;    Blue = 8'hda;
end 13'h1b:    begin Red = 8'h8b;    Green = 8'hd1;    Blue = 8'hdc;
end 13'h1c:    begin Red = 8'h91;    Green = 8'hce;    Blue = 8'he7;
end 13'h1d:    begin Red = 8'h8b;    Green = 8'hcd;    Blue = 8'hd9;
end 13'h1e:    begin Red = 8'h91;    Green = 8'hdc;    Blue = 8'hf0;
end 13'h1f:    begin Red = 8'h78;    Green = 8'h8e;    Blue = 8'h90;
end 13'h20:    begin Red = 8'h51;    Green = 8'h69;    Blue = 8'h70;
end 13'h21:    begin Red = 8'h51;    Green = 8'h5c;    Blue = 8'h5c;
end 13'h22:    begin Red = 8'h52;    Green = 8'h54;    Blue = 8'h5d;
end 13'h23:    begin Red = 8'h48;    Green = 8'h57;    Blue = 8'h5a;
end 13'h24:    begin Red = 8'h93;    Green = 8'hce;    Blue = 8'he1;
end 13'h25:    begin Red = 8'h94;    Green = 8'hc9;    Blue = 8'he5;
end 13'h26:    begin Red = 8'h7d;    Green = 8'h7f;    Blue = 8'h76;
end 13'h27:    begin Red = 8'h7d;    Green = 8'h88;    Blue = 8'h89;
end 13'h28:    begin Red = 8'h84;    Green = 8'h98;    Blue = 8'h9d;
end 13'h29:    begin Red = 8'h7c;    Green = 8'h9b;    Blue = 8'h97;
end 13'h2a:    begin Red = 8'h7a;    Green = 8'h90;    Blue = 8'h93;
end 13'h2b:    begin Red = 8'h57;    Green = 8'h6c;    Blue = 8'h72;
end 13'h2c:    begin Red = 8'h56;    Green = 8'h71;    Blue = 8'h71;
end 13'h2d:    begin Red = 8'h59;    Green = 8'h6f;    Blue = 8'h7a;
end 13'h2e:    begin Red = 8'h5f;    Green = 8'h6c;    Blue = 8'h79;
end 13'h2f:    begin Red = 8'h55;    Green = 8'h6d;    Blue = 8'h6d;
end 13'h30:    begin Red = 8'h92;    Green = 8'hca;    Blue = 8'he1;
end 13'h31:    begin Red = 8'h90;    Green = 8'hcd;    Blue = 8'hd9;
end 13'h32:    begin Red = 8'h7a;    Green = 8'h8b;    Blue = 8'h8c;
end 13'h33:    begin Red = 8'h5c;    Green = 8'h72;    Blue = 8'h75;
end 13'h34:    begin Red = 8'h61;    Green = 8'h74;    Blue = 8'h7c;
end 13'h35:    begin Red = 8'h94;    Green = 8'hdd;    Blue = 8'hf2;
end 13'h36:    begin Red = 8'h8e;    Green = 8'hc8;    Blue = 8'he2;
end 13'h37:    begin Red = 8'h90;    Green = 8'hc7;    Blue = 8'hde;
end 13'h38:    begin Red = 8'h7e;    Green = 8'h94;    Blue = 8'h9d;
end 13'h39:    begin Red = 8'h7d;    Green = 8'h98;    Blue = 8'h9a;
end 13'h3a:    begin Red = 8'h82;    Green = 8'h94;    Blue = 8'h9f;
end 13'h3b:    begin Red = 8'h5f;    Green = 8'h76;    Blue = 8'h7d;
end 13'h3c:    begin Red = 8'h63;    Green = 8'h7b;    Blue = 8'h7d;
end 13'h3d:    begin Red = 8'h58;    Green = 8'h65;    Blue = 8'h65;
end 13'h3e:    begin Red = 8'h5f;    Green = 8'h70;    Blue = 8'h71;
end 13'h3f:    begin Red = 8'h4f;    Green = 8'h6f;    Blue = 8'h6e;
end 13'h40:    begin Red = 8'h5b;    Green = 8'h69;    Blue = 8'h75;
end 13'h41:    begin Red = 8'h53;    Green = 8'h59;    Blue = 8'h5d;
end 13'h42:    begin Red = 8'h89;    Green = 8'hcd;    Blue = 8'hde;
end 13'h43:    begin Red = 8'h81;    Green = 8'h8e;    Blue = 8'h8e;
end 13'h44:    begin Red = 8'h7e;    Green = 8'h8b;    Blue = 8'h88;
end 13'h45:    begin Red = 8'h80;    Green = 8'h95;    Blue = 8'h9b;
end 13'h46:    begin Red = 8'h80;    Green = 8'h9c;    Blue = 8'h99;
end 13'h47:    begin Red = 8'h81;    Green = 8'h9a;    Blue = 8'h96;
end 13'h48:    begin Red = 8'ha6;    Green = 8'hbf;    Blue = 8'h9f;
end 13'h49:    begin Red = 8'ha3;    Green = 8'hbd;    Blue = 8'h9b;
end 13'h4a:    begin Red = 8'ha7;    Green = 8'hc1;    Blue = 8'h9b;
end 13'h4b:    begin Red = 8'h5e;    Green = 8'h75;    Blue = 8'h7a;
end 13'h4c:    begin Red = 8'h61;    Green = 8'h77;    Blue = 8'h84;
end 13'h4d:    begin Red = 8'h69;    Green = 8'h7f;    Blue = 8'h86;
end 13'h4e:    begin Red = 8'h68;    Green = 8'h7c;    Blue = 8'h81;
end 13'h4f:    begin Red = 8'h68;    Green = 8'h82;    Blue = 8'h89;
end 13'h50:    begin Red = 8'h95;    Green = 8'he4;    Blue = 8'hf6;
end 13'h51:    begin Red = 8'h92;    Green = 8'hcd;    Blue = 8'hd6;
end 13'h52:    begin Red = 8'h9a;    Green = 8'hb3;    Blue = 8'h96;
end 13'h53:    begin Red = 8'h9c;    Green = 8'hb5;    Blue = 8'h9a;
end 13'h54:    begin Red = 8'h76;    Green = 8'h8c;    Blue = 8'h8f;
end 13'h55:    begin Red = 8'h50;    Green = 8'h66;    Blue = 8'h69;
end 13'h56:    begin Red = 8'h56;    Green = 8'h5d;    Blue = 8'h65;
end 13'h57:    begin Red = 8'h4c;    Green = 8'h5b;    Blue = 8'h58;
end 13'h58:    begin Red = 8'h4b;    Green = 8'h46;    Blue = 8'h50;
end 13'h59:    begin Red = 8'h80;    Green = 8'h81;    Blue = 8'h7d;
end 13'h5a:    begin Red = 8'h79;    Green = 8'h89;    Blue = 8'h88;
end 13'h5b:    begin Red = 8'h80;    Green = 8'h93;    Blue = 8'h96;
end 13'h5c:    begin Red = 8'h83;    Green = 8'h96;    Blue = 8'h98;
end 13'h5d:    begin Red = 8'ha1;    Green = 8'hbc;    Blue = 8'h94;
end 13'h5e:    begin Red = 8'h9f;    Green = 8'hb7;    Blue = 8'h9a;
end 13'h5f:    begin Red = 8'ha6;    Green = 8'hbb;    Blue = 8'h9d;
end 13'h60:    begin Red = 8'h82;    Green = 8'h93;    Blue = 8'h7a;
end 13'h61:    begin Red = 8'h84;    Green = 8'h94;    Blue = 8'h7c;
end 13'h62:    begin Red = 8'h4f;    Green = 8'h5e;    Blue = 8'h63;
end 13'h63:    begin Red = 8'h55;    Green = 8'h75;    Blue = 8'h76;
end 13'h64:    begin Red = 8'h4e;    Green = 8'h5a;    Blue = 8'h69;
end 13'h65:    begin Red = 8'h99;    Green = 8'he5;    Blue = 8'hfd;
end 13'h66:    begin Red = 8'h89;    Green = 8'h91;    Blue = 8'h99;
end 13'h67:    begin Red = 8'h87;    Green = 8'h9e;    Blue = 8'ha1;
end 13'h68:    begin Red = 8'h80;    Green = 8'h97;    Blue = 8'ha0;
end 13'h69:    begin Red = 8'h79;    Green = 8'h91;    Blue = 8'h9a;
end 13'h6a:    begin Red = 8'h7b;    Green = 8'h90;    Blue = 8'h9e;
end 13'h6b:    begin Red = 8'h9d;    Green = 8'hbb;    Blue = 8'h91;
end 13'h6c:    begin Red = 8'h7c;    Green = 8'h8f;    Blue = 8'h7a;
end 13'h6d:    begin Red = 8'h7e;    Green = 8'h9b;    Blue = 8'h93;
end 13'h6e:    begin Red = 8'h7b;    Green = 8'h92;    Blue = 8'h95;
end 13'h6f:    begin Red = 8'h4d;    Green = 8'h5d;    Blue = 8'h60;
end 13'h70:    begin Red = 8'h4e;    Green = 8'h62;    Blue = 8'h66;
end 13'h71:    begin Red = 8'h53;    Green = 8'h63;    Blue = 8'h6a;
end 13'h72:    begin Red = 8'h56;    Green = 8'h68;    Blue = 8'h73;
end 13'h73:    begin Red = 8'h5a;    Green = 8'h71;    Blue = 8'h6d;
end 13'h74:    begin Red = 8'ha1;    Green = 8'hbd;    Blue = 8'ha3;
end 13'h75:    begin Red = 8'h99;    Green = 8'hb5;    Blue = 8'h94;
end 13'h76:    begin Red = 8'h9b;    Green = 8'hb4;    Blue = 8'h91;
end 13'h77:    begin Red = 8'ha0;    Green = 8'hb7;    Blue = 8'h9e;
end 13'h78:    begin Red = 8'ha6;    Green = 8'hbd;    Blue = 8'ha4;
end 13'h79:    begin Red = 8'h82;    Green = 8'h94;    Blue = 8'h80;
end 13'h7a:    begin Red = 8'h83;    Green = 8'h95;    Blue = 8'ha2;
end 13'h7b:    begin Red = 8'h62;    Green = 8'h7a;    Blue = 8'h83;
end 13'h7c:    begin Red = 8'h62;    Green = 8'h79;    Blue = 8'h88;
end 13'h7d:    begin Red = 8'h6c;    Green = 8'h80;    Blue = 8'h84;
end 13'h7e:    begin Red = 8'h5e;    Green = 8'h70;    Blue = 8'h78;
end 13'h7f:    begin Red = 8'h5e;    Green = 8'h6e;    Blue = 8'h74;
end 13'h80:    begin Red = 8'h5c;    Green = 8'h6d;    Blue = 8'h76;
end 13'h81:    begin Red = 8'h4a;    Green = 8'h61;    Blue = 8'h64;
end 13'h82:    begin Red = 8'h7d;    Green = 8'h96;    Blue = 8'h91;
end 13'h83:    begin Red = 8'h9d;    Green = 8'hb3;    Blue = 8'h93;
end 13'h84:    begin Red = 8'h9b;    Green = 8'hb2;    Blue = 8'h9b;
end 13'h85:    begin Red = 8'h9d;    Green = 8'hb5;    Blue = 8'h9f;
end 13'h86:    begin Red = 8'ha3;    Green = 8'hbb;    Blue = 8'h9f;
end 13'h87:    begin Red = 8'hac;    Green = 8'hbf;    Blue = 8'ha7;
end 13'h88:    begin Red = 8'h81;    Green = 8'h91;    Blue = 8'h7d;
end 13'h89:    begin Red = 8'h83;    Green = 8'h99;    Blue = 8'h79;
end 13'h8a:    begin Red = 8'h85;    Green = 8'h97;    Blue = 8'h78;
end 13'h8b:    begin Red = 8'h66;    Green = 8'h79;    Blue = 8'h7d;
end 13'h8c:    begin Red = 8'h6a;    Green = 8'h78;    Blue = 8'h82;
end 13'h8d:    begin Red = 8'hdc;    Green = 8'hd9;    Blue = 8'hce;
end 13'h8e:    begin Red = 8'hca;    Green = 8'hc7;    Blue = 8'hbb;
end 13'h8f:    begin Red = 8'hca;    Green = 8'hc3;    Blue = 8'hb9;
end 13'h90:    begin Red = 8'hd4;    Green = 8'hce;    Blue = 8'hc3;
end 13'h91:    begin Red = 8'hcf;    Green = 8'hca;    Blue = 8'hbf;
end 13'h92:    begin Red = 8'h52;    Green = 8'h69;    Blue = 8'h6c;
end 13'h93:    begin Red = 8'h9c;    Green = 8'hb7;    Blue = 8'h94;
end 13'h94:    begin Red = 8'h65;    Green = 8'h78;    Blue = 8'h86;
end 13'h95:    begin Red = 8'h66;    Green = 8'h79;    Blue = 8'h83;
end 13'h96:    begin Red = 8'h65;    Green = 8'h7c;    Blue = 8'h7a;
end 13'h97:    begin Red = 8'hc7;    Green = 8'hc7;    Blue = 8'hbf;
end 13'h98:    begin Red = 8'hca;    Green = 8'hca;    Blue = 8'hc2;
end 13'h99:    begin Red = 8'hb8;    Green = 8'hb8;    Blue = 8'hb0;
end 13'h9a:    begin Red = 8'h9c;    Green = 8'hb3;    Blue = 8'ha2;
end 13'h9b:    begin Red = 8'h87;    Green = 8'h94;    Blue = 8'h7f;
end 13'h9c:    begin Red = 8'h83;    Green = 8'h97;    Blue = 8'h7d;
end 13'h9d:    begin Red = 8'hc5;    Green = 8'hca;    Blue = 8'hbe;
end 13'h9e:    begin Red = 8'hc3;    Green = 8'hc7;    Blue = 8'hc4;
end 13'h9f:    begin Red = 8'h7a;    Green = 8'h8d;    Blue = 8'h7c;
end 13'ha0:    begin Red = 8'h79;    Green = 8'h8e;    Blue = 8'h77;
end 13'ha1:    begin Red = 8'h7d;    Green = 8'h97;    Blue = 8'h9e;
end 13'ha2:    begin Red = 8'h5d;    Green = 8'h76;    Blue = 8'h82;
end 13'ha3:    begin Red = 8'h63;    Green = 8'h7f;    Blue = 8'h84;
end 13'ha4:    begin Red = 8'h4a;    Green = 8'h6c;    Blue = 8'h75;
end 13'ha5:    begin Red = 8'h50;    Green = 8'h6d;    Blue = 8'h82;
end 13'ha6:    begin Red = 8'h51;    Green = 8'h6a;    Blue = 8'h76;
end 13'ha7:    begin Red = 8'hc6;    Green = 8'hc8;    Blue = 8'hc3;
end 13'ha8:    begin Red = 8'hbd;    Green = 8'hc3;    Blue = 8'hbd;
end 13'ha9:    begin Red = 8'hba;    Green = 8'hc5;    Blue = 8'hb7;
end 13'haa:    begin Red = 8'h88;    Green = 8'ha1;    Blue = 8'ha3;
end 13'hab:    begin Red = 8'h7e;    Green = 8'h98;    Blue = 8'h8f;
end 13'hac:    begin Red = 8'h8e;    Green = 8'h9b;    Blue = 8'h77;
end 13'had:    begin Red = 8'h64;    Green = 8'h7b;    Blue = 8'h89;
end 13'hae:    begin Red = 8'h55;    Green = 8'h7a;    Blue = 8'h78;
end 13'haf:    begin Red = 8'ha7;    Green = 8'h8d;    Blue = 8'h75;
end 13'hb0:    begin Red = 8'hbb;    Green = 8'hba;    Blue = 8'hb7;
end 13'hb1:    begin Red = 8'hb5;    Green = 8'hb9;    Blue = 8'hb6;
end 13'hb2:    begin Red = 8'ha0;    Green = 8'h86;    Blue = 8'h65;
end 13'hb3:    begin Red = 8'ha4;    Green = 8'haf;    Blue = 8'ha7;
end 13'hb4:    begin Red = 8'ha6;    Green = 8'ha0;    Blue = 8'h91;
end 13'hb5:    begin Red = 8'hb7;    Green = 8'hbc;    Blue = 8'hb4;
end 13'hb6:    begin Red = 8'hba;    Green = 8'hba;    Blue = 8'hb2;
end 13'hb7:    begin Red = 8'hb5;    Green = 8'hb5;    Blue = 8'had;
end 13'hb8:    begin Red = 8'h7b;    Green = 8'h8c;    Blue = 8'h83;
end 13'hb9:    begin Red = 8'h84;    Green = 8'h95;    Blue = 8'h83;
end 13'hba:    begin Red = 8'h80;    Green = 8'h94;    Blue = 8'h85;
end 13'hbb:    begin Red = 8'h60;    Green = 8'h72;    Blue = 8'h77;
end 13'hbc:    begin Red = 8'h5e;    Green = 8'h71;    Blue = 8'h7c;
end 13'hbd:    begin Red = 8'hb7;    Green = 8'h99;    Blue = 8'h74;
end 13'hbe:    begin Red = 8'hb9;    Green = 8'h9d;    Blue = 8'h7c;
end 13'hbf:    begin Red = 8'hac;    Green = 8'h8f;    Blue = 8'h72;
end 13'hc0:    begin Red = 8'hbf;    Green = 8'hb9;    Blue = 8'hb7;
end 13'hc1:    begin Red = 8'hcc;    Green = 8'hcc;    Blue = 8'hc4;
end 13'hc2:    begin Red = 8'h98;    Green = 8'h84;    Blue = 8'h6e;
end 13'hc3:    begin Red = 8'ha3;    Green = 8'h90;    Blue = 8'h70;
end 13'hc4:    begin Red = 8'haa;    Green = 8'ha5;    Blue = 8'h9b;
end 13'hc5:    begin Red = 8'ha0;    Green = 8'ha0;    Blue = 8'h98;
end 13'hc6:    begin Red = 8'h5c;    Green = 8'h70;    Blue = 8'h80;
end 13'hc7:    begin Red = 8'hba;    Green = 8'h9a;    Blue = 8'h73;
end 13'hc8:    begin Red = 8'hbe;    Green = 8'h9a;    Blue = 8'h7d;
end 13'hc9:    begin Red = 8'h9b;    Green = 8'h84;    Blue = 8'h69;
end 13'hca:    begin Red = 8'haf;    Green = 8'h8c;    Blue = 8'h75;
end 13'hcb:    begin Red = 8'ha4;    Green = 8'h90;    Blue = 8'h78;
end 13'hcc:    begin Red = 8'ha4;    Green = 8'ha7;    Blue = 8'h99;
end 13'hcd:    begin Red = 8'ha1;    Green = 8'h9e;    Blue = 8'h8a;
end 13'hce:    begin Red = 8'hbe;    Green = 8'hb6;    Blue = 8'hb1;
end 13'hcf:    begin Red = 8'h98;    Green = 8'hb1;    Blue = 8'h9f;
end 13'hd0:    begin Red = 8'hce;    Green = 8'h9e;    Blue = 8'h7b;
end 13'hd1:    begin Red = 8'hbb;    Green = 8'h98;    Blue = 8'h7d;
end 13'hd2:    begin Red = 8'ha9;    Green = 8'h8a;    Blue = 8'h68;
end 13'hd3:    begin Red = 8'ha7;    Green = 8'h8b;    Blue = 8'h71;
end 13'hd4:    begin Red = 8'ha7;    Green = 8'h89;    Blue = 8'h74;
end 13'hd5:    begin Red = 8'ha2;    Green = 8'ha2;    Blue = 8'h9a;
end 13'hd6:    begin Red = 8'hb2;    Green = 8'hba;    Blue = 8'hb1;
end 13'hd7:    begin Red = 8'h41;    Green = 8'h65;    Blue = 8'h71;
end 13'hd8:    begin Red = 8'hc5;    Green = 8'haa;    Blue = 8'h8c;
end 13'hd9:    begin Red = 8'hca;    Green = 8'hac;    Blue = 8'h8d;
end 13'hda:    begin Red = 8'h75;    Green = 8'h98;    Blue = 8'h99;
end 13'hdb:    begin Red = 8'h84;    Green = 8'h94;    Blue = 8'h95;
end 13'hdc:    begin Red = 8'h80;    Green = 8'h94;    Blue = 8'h92;
end 13'hdd:    begin Red = 8'h72;    Green = 8'h8a;    Blue = 8'h8c;
end 13'hde:    begin Red = 8'h78;    Green = 8'h8b;    Blue = 8'h93;
end 13'hdf:    begin Red = 8'had;    Green = 8'hca;    Blue = 8'h92;
end 13'he0:    begin Red = 8'h84;    Green = 8'h98;    Blue = 8'h80;
end 13'he1:    begin Red = 8'h8c;    Green = 8'h9b;    Blue = 8'h82;
end 13'he2:    begin Red = 8'h90;    Green = 8'ha0;    Blue = 8'h7b;
end 13'he3:    begin Red = 8'h61;    Green = 8'h79;    Blue = 8'h7b;
end 13'he4:    begin Red = 8'hc2;    Green = 8'h9b;    Blue = 8'h7f;
end 13'he5:    begin Red = 8'haa;    Green = 8'h8e;    Blue = 8'h76;
end 13'he6:    begin Red = 8'ha8;    Green = 8'ha8;    Blue = 8'ha0;
end 13'he7:    begin Red = 8'hb5;    Green = 8'hb6;    Blue = 8'ha9;
end 13'he8:    begin Red = 8'hac;    Green = 8'h88;    Blue = 8'h69;
end 13'he9:    begin Red = 8'h93;    Green = 8'h93;    Blue = 8'h89;
end 13'hea:    begin Red = 8'ha7;    Green = 8'ha7;    Blue = 8'h9d;
end 13'heb:    begin Red = 8'h45;    Green = 8'h61;    Blue = 8'h6b;
end 13'hec:    begin Red = 8'hbb;    Green = 8'ha4;    Blue = 8'h8b;
end 13'hed:    begin Red = 8'hbb;    Green = 8'ha7;    Blue = 8'h8f;
end 13'hee:    begin Red = 8'h7e;    Green = 8'h9a;    Blue = 8'h9f;
end 13'hef:    begin Red = 8'ha1;    Green = 8'hba;    Blue = 8'h97;
end 13'hf0:    begin Red = 8'h88;    Green = 8'h98;    Blue = 8'h82;
end 13'hf1:    begin Red = 8'h5c;    Green = 8'h72;    Blue = 8'h85;
end 13'hf2:    begin Red = 8'hcb;    Green = 8'h9f;    Blue = 8'h78;
end 13'hf3:    begin Red = 8'haf;    Green = 8'haf;    Blue = 8'ha7;
end 13'hf4:    begin Red = 8'hac;    Green = 8'hac;    Blue = 8'ha3;
end 13'hf5:    begin Red = 8'haf;    Green = 8'h8c;    Blue = 8'h6b;
end 13'hf6:    begin Red = 8'h99;    Green = 8'h98;    Blue = 8'h8e;
end 13'hf7:    begin Red = 8'haa;    Green = 8'hab;    Blue = 8'h9e;
end 13'hf8:    begin Red = 8'ha7;    Green = 8'h94;    Blue = 8'h79;
end 13'hf9:    begin Red = 8'hb4;    Green = 8'haf;    Blue = 8'h98;
end 13'hfa:    begin Red = 8'hc1;    Green = 8'ha7;    Blue = 8'h86;
end 13'hfb:    begin Red = 8'hbc;    Green = 8'ha7;    Blue = 8'h94;
end 13'hfc:    begin Red = 8'hb7;    Green = 8'ha7;    Blue = 8'h94;
end 13'hfd:    begin Red = 8'hbe;    Green = 8'haa;    Blue = 8'h8e;
end 13'hfe:    begin Red = 8'ha3;    Green = 8'h98;    Blue = 8'h83;
end 13'hff:    begin Red = 8'h78;    Green = 8'h8e;    Blue = 8'h95;
end 13'h100:    begin Red = 8'ha4;    Green = 8'hc0;    Blue = 8'h94;
end 13'h101:    begin Red = 8'h9b;    Green = 8'hb7;    Blue = 8'h9c;
end 13'h102:    begin Red = 8'h83;    Green = 8'h95;    Blue = 8'h88;
end 13'h103:    begin Red = 8'h80;    Green = 8'h98;    Blue = 8'h84;
end 13'h104:    begin Red = 8'h88;    Green = 8'h9d;    Blue = 8'h7d;
end 13'h105:    begin Red = 8'hb7;    Green = 8'h98;    Blue = 8'h79;
end 13'h106:    begin Red = 8'hbc;    Green = 8'h98;    Blue = 8'h79;
end 13'h107:    begin Red = 8'h9a;    Green = 8'h81;    Blue = 8'h6a;
end 13'h108:    begin Red = 8'haa;    Green = 8'h88;    Blue = 8'h66;
end 13'h109:    begin Red = 8'h44;    Green = 8'h62;    Blue = 8'h71;
end 13'h10a:    begin Red = 8'h39;    Green = 8'h5e;    Blue = 8'h75;
end 13'h10b:    begin Red = 8'ha7;    Green = 8'h99;    Blue = 8'h86;
end 13'h10c:    begin Red = 8'hbf;    Green = 8'hac;    Blue = 8'h93;
end 13'h10d:    begin Red = 8'hbb;    Green = 8'ha8;    Blue = 8'h8a;
end 13'h10e:    begin Red = 8'ha6;    Green = 8'h95;    Blue = 8'h80;
end 13'h10f:    begin Red = 8'h71;    Green = 8'h92;    Blue = 8'h9d;
end 13'h110:    begin Red = 8'h6d;    Green = 8'h92;    Blue = 8'h9f;
end 13'h111:    begin Red = 8'h77;    Green = 8'h8f;    Blue = 8'h88;
end 13'h112:    begin Red = 8'h71;    Green = 8'h86;    Blue = 8'h8c;
end 13'h113:    begin Red = 8'h89;    Green = 8'h9f;    Blue = 8'h83;
end 13'h114:    begin Red = 8'h5e;    Green = 8'h74;    Blue = 8'h84;
end 13'h115:    begin Red = 8'h5a;    Green = 8'h74;    Blue = 8'h80;
end 13'h116:    begin Red = 8'hbb;    Green = 8'h9b;    Blue = 8'h7b;
end 13'h117:    begin Red = 8'ha7;    Green = 8'h84;    Blue = 8'h63;
end 13'h118:    begin Red = 8'hbe;    Green = 8'hbe;    Blue = 8'hb6;
end 13'h119:    begin Red = 8'ha4;    Green = 8'h94;    Blue = 8'h7e;
end 13'h11a:    begin Red = 8'hbf;    Green = 8'ha7;    Blue = 8'h90;
end 13'h11b:    begin Red = 8'h77;    Green = 8'h90;    Blue = 8'h8c;
end 13'h11c:    begin Red = 8'h71;    Green = 8'h87;    Blue = 8'h90;
end 13'h11d:    begin Red = 8'h86;    Green = 8'h98;    Blue = 8'h85;
end 13'h11e:    begin Red = 8'h8a;    Green = 8'h9a;    Blue = 8'h7d;
end 13'h11f:    begin Red = 8'h9f;    Green = 8'h9f;    Blue = 8'h95;
end 13'h120:    begin Red = 8'h59;    Green = 8'h74;    Blue = 8'h75;
end 13'h121:    begin Red = 8'h78;    Green = 8'h96;    Blue = 8'h98;
end 13'h122:    begin Red = 8'h86;    Green = 8'h98;    Blue = 8'ha3;
end 13'h123:    begin Red = 8'h7b;    Green = 8'h90;    Blue = 8'ha3;
end 13'h124:    begin Red = 8'h61;    Green = 8'h7e;    Blue = 8'h73;
end 13'h125:    begin Red = 8'hf6;    Green = 8'hf0;    Blue = 8'hc4;
end 13'h126:    begin Red = 8'he2;    Green = 8'hde;    Blue = 8'hbe;
end 13'h127:    begin Red = 8'he1;    Green = 8'he2;    Blue = 8'hc3;
end 13'h128:    begin Red = 8'ha0;    Green = 8'ha7;    Blue = 8'h9a;
end 13'h129:    begin Red = 8'ha5;    Green = 8'hac;    Blue = 8'h9d;
end 13'h12a:    begin Red = 8'h93;    Green = 8'h99;    Blue = 8'h8d;
end 13'h12b:    begin Red = 8'h90;    Green = 8'h9f;    Blue = 8'h92;
end 13'h12c:    begin Red = 8'h95;    Green = 8'h9f;    Blue = 8'h94;
end 13'h12d:    begin Red = 8'hb8;    Green = 8'hbb;    Blue = 8'haa;
end 13'h12e:    begin Red = 8'h98;    Green = 8'h9a;    Blue = 8'h89;
end 13'h12f:    begin Red = 8'h8a;    Green = 8'h95;    Blue = 8'h81;
end 13'h130:    begin Red = 8'h8f;    Green = 8'h98;    Blue = 8'h8a;
end 13'h131:    begin Red = 8'h90;    Green = 8'h98;    Blue = 8'h84;
end 13'h132:    begin Red = 8'h8a;    Green = 8'h8a;    Blue = 8'h82;
end 13'h133:    begin Red = 8'h8c;    Green = 8'h82;    Blue = 8'h7b;
end 13'h134:    begin Red = 8'h80;    Green = 8'h83;    Blue = 8'h6f;
end 13'h135:    begin Red = 8'h4b;    Green = 8'h6b;    Blue = 8'h71;
end 13'h136:    begin Red = 8'h35;    Green = 8'h57;    Blue = 8'h66;
end 13'h137:    begin Red = 8'h3a;    Green = 8'h55;    Blue = 8'h62;
end 13'h138:    begin Red = 8'h71;    Green = 8'h8c;    Blue = 8'h93;
end 13'h139:    begin Red = 8'h5e;    Green = 8'h85;    Blue = 8'h90;
end 13'h13a:    begin Red = 8'h61;    Green = 8'h88;    Blue = 8'h95;
end 13'h13b:    begin Red = 8'h65;    Green = 8'h87;    Blue = 8'h90;
end 13'h13c:    begin Red = 8'h67;    Green = 8'h85;    Blue = 8'h8c;
end 13'h13d:    begin Red = 8'h6a;    Green = 8'h87;    Blue = 8'h92;
end 13'h13e:    begin Red = 8'h76;    Green = 8'h8b;    Blue = 8'h9d;
end 13'h13f:    begin Red = 8'h7f;    Green = 8'h93;    Blue = 8'h7c;
end 13'h140:    begin Red = 8'h7f;    Green = 8'h99;    Blue = 8'h77;
end 13'h141:    begin Red = 8'he8;    Green = 8'hde;    Blue = 8'hb8;
end 13'h142:    begin Red = 8'hcd;    Green = 8'hcd;    Blue = 8'hb8;
end 13'h143:    begin Red = 8'hc7;    Green = 8'hc9;    Blue = 8'hac;
end 13'h144:    begin Red = 8'h9f;    Green = 8'h9d;    Blue = 8'h8c;
end 13'h145:    begin Red = 8'ha8;    Green = 8'ha8;    Blue = 8'h92;
end 13'h146:    begin Red = 8'h95;    Green = 8'h9e;    Blue = 8'h84;
end 13'h147:    begin Red = 8'h9b;    Green = 8'h98;    Blue = 8'h88;
end 13'h148:    begin Red = 8'h98;    Green = 8'h90;    Blue = 8'h80;
end 13'h149:    begin Red = 8'h94;    Green = 8'h94;    Blue = 8'h84;
end 13'h14a:    begin Red = 8'ha1;    Green = 8'h91;    Blue = 8'h8c;
end 13'h14b:    begin Red = 8'h86;    Green = 8'h88;    Blue = 8'h7d;
end 13'h14c:    begin Red = 8'h88;    Green = 8'h8c;    Blue = 8'h80;
end 13'h14d:    begin Red = 8'h86;    Green = 8'h86;    Blue = 8'h73;
end 13'h14e:    begin Red = 8'h61;    Green = 8'h7b;    Blue = 8'h8d;
end 13'h14f:    begin Red = 8'h65;    Green = 8'h7d;    Blue = 8'h7e;
end 13'h150:    begin Red = 8'h5e;    Green = 8'h6c;    Blue = 8'h6e;
end 13'h151:    begin Red = 8'h61;    Green = 8'h6f;    Blue = 8'h75;
end 13'h152:    begin Red = 8'hf3;    Green = 8'hde;    Blue = 8'hbb;
end 13'h153:    begin Red = 8'h55;    Green = 8'h70;    Blue = 8'h74;
end 13'h154:    begin Red = 8'hc2;    Green = 8'haa;    Blue = 8'h97;
end 13'h155:    begin Red = 8'hc7;    Green = 8'hac;    Blue = 8'h88;
end 13'h156:    begin Red = 8'hfb;    Green = 8'hed;    Blue = 8'hc4;
end 13'h157:    begin Red = 8'hf1;    Green = 8'hde;    Blue = 8'hbf;
end 13'h158:    begin Red = 8'hf1;    Green = 8'he0;    Blue = 8'hbc;
end 13'h159:    begin Red = 8'ha0;    Green = 8'hb3;    Blue = 8'h9a;
end 13'h15a:    begin Red = 8'h99;    Green = 8'hb6;    Blue = 8'h99;
end 13'h15b:    begin Red = 8'ha0;    Green = 8'hb3;    Blue = 8'ha0;
end 13'h15c:    begin Red = 8'ha4;    Green = 8'hbb;    Blue = 8'ha3;
end 13'h15d:    begin Red = 8'h60;    Green = 8'h80;    Blue = 8'h79;
end 13'h15e:    begin Red = 8'he0;    Green = 8'hdd;    Blue = 8'hb9;
end 13'h15f:    begin Red = 8'hca;    Green = 8'hca;    Blue = 8'hab;
end 13'h160:    begin Red = 8'ha6;    Green = 8'ha5;    Blue = 8'h95;
end 13'h161:    begin Red = 8'h9b;    Green = 8'h9b;    Blue = 8'h8b;
end 13'h162:    begin Red = 8'hc4;    Green = 8'hc4;    Blue = 8'hbc;
end 13'h163:    begin Red = 8'h98;    Green = 8'h97;    Blue = 8'h87;
end 13'h164:    begin Red = 8'h8c;    Green = 8'h8a;    Blue = 8'h7e;
end 13'h165:    begin Red = 8'h87;    Green = 8'h85;    Blue = 8'h79;
end 13'h166:    begin Red = 8'h61;    Green = 8'h6f;    Blue = 8'h8d;
end 13'h167:    begin Red = 8'ha6;    Green = 8'hb7;    Blue = 8'h56;
end 13'h168:    begin Red = 8'ha5;    Green = 8'hb3;    Blue = 8'h54;
end 13'h169:    begin Red = 8'hfe;    Green = 8'hff;    Blue = 8'hd9;
end 13'h16a:    begin Red = 8'hff;    Green = 8'hf9;    Blue = 8'hcb;
end 13'h16b:    begin Red = 8'hff;    Green = 8'hf4;    Blue = 8'hd6;
end 13'h16c:    begin Red = 8'hfa;    Green = 8'hf1;    Blue = 8'hc3;
end 13'h16d:    begin Red = 8'hf2;    Green = 8'he2;    Blue = 8'hbe;
end 13'h16e:    begin Red = 8'hf8;    Green = 8'hd9;    Blue = 8'hac;
end 13'h16f:    begin Red = 8'hf6;    Green = 8'hd9;    Blue = 8'hb3;
end 13'h170:    begin Red = 8'hff;    Green = 8'hf5;    Blue = 8'hca;
end 13'h171:    begin Red = 8'hff;    Green = 8'hfb;    Blue = 8'hce;
end 13'h172:    begin Red = 8'hb3;    Green = 8'hac;    Blue = 8'h8c;
end 13'h173:    begin Red = 8'ha3;    Green = 8'h8f;    Blue = 8'h75;
end 13'h174:    begin Red = 8'h7a;    Green = 8'h67;    Blue = 8'h51;
end 13'h175:    begin Red = 8'h80;    Green = 8'h6f;    Blue = 8'h5a;
end 13'h176:    begin Red = 8'h7e;    Green = 8'h6c;    Blue = 8'h53;
end 13'h177:    begin Red = 8'hb9;    Green = 8'ha3;    Blue = 8'h92;
end 13'h178:    begin Red = 8'hf0;    Green = 8'hcd;    Blue = 8'ha7;
end 13'h179:    begin Red = 8'hf5;    Green = 8'hf5;    Blue = 8'hcb;
end 13'h17a:    begin Red = 8'hff;    Green = 8'hed;    Blue = 8'hc5;
end 13'h17b:    begin Red = 8'hff;    Green = 8'hdb;    Blue = 8'hbb;
end 13'h17c:    begin Red = 8'hf6;    Green = 8'hdf;    Blue = 8'hbe;
end 13'h17d:    begin Red = 8'hee;    Green = 8'hde;    Blue = 8'hc7;
end 13'h17e:    begin Red = 8'hf1;    Green = 8'hdc;    Blue = 8'hb8;
end 13'h17f:    begin Red = 8'hff;    Green = 8'he6;    Blue = 8'hc1;
end 13'h180:    begin Red = 8'h95;    Green = 8'ha9;    Blue = 8'h91;
end 13'h181:    begin Red = 8'hfd;    Green = 8'hf8;    Blue = 8'hf8;
end 13'h182:    begin Red = 8'hf9;    Green = 8'hf2;    Blue = 8'hf6;
end 13'h183:    begin Red = 8'hfc;    Green = 8'hf4;    Blue = 8'hfa;
end 13'h184:    begin Red = 8'hff;    Green = 8'hfc;    Blue = 8'hff;
end 13'h185:    begin Red = 8'hfd;    Green = 8'hfd;    Blue = 8'hfd;
end 13'h186:    begin Red = 8'hf9;    Green = 8'hf5;    Blue = 8'hf8;
end 13'h187:    begin Red = 8'h77;    Green = 8'h8c;    Blue = 8'h76;
end 13'h188:    begin Red = 8'h8d;    Green = 8'haa;    Blue = 8'h8d;
end 13'h189:    begin Red = 8'h80;    Green = 8'h8e;    Blue = 8'h81;
end 13'h18a:    begin Red = 8'h7d;    Green = 8'h90;    Blue = 8'h7f;
end 13'h18b:    begin Red = 8'h53;    Green = 8'h74;    Blue = 8'h8d;
end 13'h18c:    begin Red = 8'h9a;    Green = 8'ha7;    Blue = 8'h60;
end 13'h18d:    begin Red = 8'h97;    Green = 8'ha7;    Blue = 8'h5c;
end 13'h18e:    begin Red = 8'h96;    Green = 8'ha6;    Blue = 8'h5f;
end 13'h18f:    begin Red = 8'hff;    Green = 8'hf6;    Blue = 8'hd2;
end 13'h190:    begin Red = 8'hf7;    Green = 8'hdb;    Blue = 8'hbb;
end 13'h191:    begin Red = 8'hf1;    Green = 8'hde;    Blue = 8'hac;
end 13'h192:    begin Red = 8'hd8;    Green = 8'hc4;    Blue = 8'ha4;
end 13'h193:    begin Red = 8'hda;    Green = 8'hc3;    Blue = 8'ha6;
end 13'h194:    begin Red = 8'hf1;    Green = 8'hdd;    Blue = 8'hc4;
end 13'h195:    begin Red = 8'hbc;    Green = 8'had;    Blue = 8'h94;
end 13'h196:    begin Red = 8'h85;    Green = 8'h74;    Blue = 8'h61;
end 13'h197:    begin Red = 8'h82;    Green = 8'h6e;    Blue = 8'h5d;
end 13'h198:    begin Red = 8'h8b;    Green = 8'h7b;    Blue = 8'h68;
end 13'h199:    begin Red = 8'hb6;    Green = 8'ha0;    Blue = 8'h90;
end 13'h19a:    begin Red = 8'hd9;    Green = 8'hc6;    Blue = 8'ha0;
end 13'h19b:    begin Red = 8'hf8;    Green = 8'he6;    Blue = 8'hc7;
end 13'h19c:    begin Red = 8'heb;    Green = 8'he2;    Blue = 8'hc3;
end 13'h19d:    begin Red = 8'hee;    Green = 8'hdf;    Blue = 8'hbe;
end 13'h19e:    begin Red = 8'ha8;    Green = 8'hb2;    Blue = 8'h9f;
end 13'h19f:    begin Red = 8'h83;    Green = 8'hae;    Blue = 8'h84;
end 13'h1a0:    begin Red = 8'hf1;    Green = 8'hea;    Blue = 8'hea;
end 13'h1a1:    begin Red = 8'heb;    Green = 8'he9;    Blue = 8'he5;
end 13'h1a2:    begin Red = 8'he7;    Green = 8'he7;    Blue = 8'he7;
end 13'h1a3:    begin Red = 8'hed;    Green = 8'hed;    Blue = 8'hea;
end 13'h1a4:    begin Red = 8'hfe;    Green = 8'hf1;    Blue = 8'hf9;
end 13'h1a5:    begin Red = 8'hfe;    Green = 8'hf3;    Blue = 8'hf3;
end 13'h1a6:    begin Red = 8'heb;    Green = 8'hec;    Blue = 8'he7;
end 13'h1a7:    begin Red = 8'he7;    Green = 8'he6;    Blue = 8'he3;
end 13'h1a8:    begin Red = 8'h80;    Green = 8'h95;    Blue = 8'h7e;
end 13'h1a9:    begin Red = 8'h8a;    Green = 8'ha8;    Blue = 8'h89;
end 13'h1aa:    begin Red = 8'h7e;    Green = 8'h97;    Blue = 8'h7d;
end 13'h1ab:    begin Red = 8'h64;    Green = 8'h7c;    Blue = 8'h8f;
end 13'h1ac:    begin Red = 8'h83;    Green = 8'h97;    Blue = 8'h55;
end 13'h1ad:    begin Red = 8'h64;    Green = 8'h7d;    Blue = 8'h76;
end 13'h1ae:    begin Red = 8'h68;    Green = 8'h7a;    Blue = 8'h88;
end 13'h1af:    begin Red = 8'h8e;    Green = 8'h99;    Blue = 8'h54;
end 13'h1b0:    begin Red = 8'h87;    Green = 8'h93;    Blue = 8'h5c;
end 13'h1b1:    begin Red = 8'h95;    Green = 8'ha7;    Blue = 8'h59;
end 13'h1b2:    begin Red = 8'h85;    Green = 8'h93;    Blue = 8'h53;
end 13'h1b3:    begin Red = 8'h71;    Green = 8'h7b;    Blue = 8'h4a;
end 13'h1b4:    begin Red = 8'h66;    Green = 8'h77;    Blue = 8'h48;
end 13'h1b5:    begin Red = 8'h99;    Green = 8'hab;    Blue = 8'h55;
end 13'h1b6:    begin Red = 8'hfd;    Green = 8'he7;    Blue = 8'hc5;
end 13'h1b7:    begin Red = 8'hf7;    Green = 8'he3;    Blue = 8'hc3;
end 13'h1b8:    begin Red = 8'hff;    Green = 8'hee;    Blue = 8'hce;
end 13'h1b9:    begin Red = 8'ha4;    Green = 8'h93;    Blue = 8'h74;
end 13'h1ba:    begin Red = 8'hcf;    Green = 8'hbe;    Blue = 8'h98;
end 13'h1bb:    begin Red = 8'hc7;    Green = 8'hb3;    Blue = 8'h93;
end 13'h1bc:    begin Red = 8'hc3;    Green = 8'hb2;    Blue = 8'h94;
end 13'h1bd:    begin Red = 8'hdd;    Green = 8'hc7;    Blue = 8'ha5;
end 13'h1be:    begin Red = 8'hf4;    Green = 8'hdf;    Blue = 8'hb8;
end 13'h1bf:    begin Red = 8'hac;    Green = 8'h98;    Blue = 8'h80;
end 13'h1c0:    begin Red = 8'h8c;    Green = 8'h7c;    Blue = 8'h65;
end 13'h1c1:    begin Red = 8'hac;    Green = 8'h96;    Blue = 8'h83;
end 13'h1c2:    begin Red = 8'ha4;    Green = 8'h8e;    Blue = 8'h7b;
end 13'h1c3:    begin Red = 8'hb5;    Green = 8'ha4;    Blue = 8'h8c;
end 13'h1c4:    begin Red = 8'hdc;    Green = 8'hcb;    Blue = 8'ha7;
end 13'h1c5:    begin Red = 8'hf7;    Green = 8'he2;    Blue = 8'hbf;
end 13'h1c6:    begin Red = 8'hb7;    Green = 8'ha4;    Blue = 8'h81;
end 13'h1c7:    begin Red = 8'hc3;    Green = 8'hb0;    Blue = 8'h8f;
end 13'h1c8:    begin Red = 8'ha1;    Green = 8'h8e;    Blue = 8'h73;
end 13'h1c9:    begin Red = 8'ha3;    Green = 8'hb7;    Blue = 8'ha0;
end 13'h1ca:    begin Red = 8'heb;    Green = 8'he8;    Blue = 8'he9;
end 13'h1cb:    begin Red = 8'hff;    Green = 8'hf9;    Blue = 8'hfd;
end 13'h1cc:    begin Red = 8'h85;    Green = 8'h91;    Blue = 8'h82;
end 13'h1cd:    begin Red = 8'h88;    Green = 8'h93;    Blue = 8'h83;
end 13'h1ce:    begin Red = 8'hea;    Green = 8'he3;    Blue = 8'he2;
end 13'h1cf:    begin Red = 8'he4;    Green = 8'hea;    Blue = 8'he0;
end 13'h1d0:    begin Red = 8'he9;    Green = 8'he9;    Blue = 8'hef;
end 13'h1d1:    begin Red = 8'hea;    Green = 8'he5;    Blue = 8'he6;
end 13'h1d2:    begin Red = 8'he4;    Green = 8'he2;    Blue = 8'he6;
end 13'h1d3:    begin Red = 8'hfb;    Green = 8'hf6;    Blue = 8'hfc;
end 13'h1d4:    begin Red = 8'h89;    Green = 8'haa;    Blue = 8'h87;
end 13'h1d5:    begin Red = 8'h86;    Green = 8'h9b;    Blue = 8'h7b;
end 13'h1d6:    begin Red = 8'h99;    Green = 8'hb0;    Blue = 8'h98;
end 13'h1d7:    begin Red = 8'h61;    Green = 8'h7d;    Blue = 8'h80;
end 13'h1d8:    begin Red = 8'hd2;    Green = 8'hd2;    Blue = 8'hb1;
end 13'h1d9:    begin Red = 8'ha4;    Green = 8'ha3;    Blue = 8'h92;
end 13'h1da:    begin Red = 8'h5d;    Green = 8'h7b;    Blue = 8'h8c;
end 13'h1db:    begin Red = 8'h56;    Green = 8'h74;    Blue = 8'h95;
end 13'h1dc:    begin Red = 8'h5a;    Green = 8'h77;    Blue = 8'h8c;
end 13'h1dd:    begin Red = 8'h5c;    Green = 8'h75;    Blue = 8'h94;
end 13'h1de:    begin Red = 8'h5c;    Green = 8'h7d;    Blue = 8'h88;
end 13'h1df:    begin Red = 8'h94;    Green = 8'ha0;    Blue = 8'h55;
end 13'h1e0:    begin Red = 8'h8e;    Green = 8'h98;    Blue = 8'h61;
end 13'h1e1:    begin Red = 8'h9a;    Green = 8'haa;    Blue = 8'h5d;
end 13'h1e2:    begin Red = 8'h85;    Green = 8'h90;    Blue = 8'h58;
end 13'h1e3:    begin Red = 8'h87;    Green = 8'h92;    Blue = 8'h55;
end 13'h1e4:    begin Red = 8'h6d;    Green = 8'h75;    Blue = 8'h4a;
end 13'h1e5:    begin Red = 8'h62;    Green = 8'h6d;    Blue = 8'h45;
end 13'h1e6:    begin Red = 8'ha0;    Green = 8'haf;    Blue = 8'h4f;
end 13'h1e7:    begin Red = 8'hfb;    Green = 8'he6;    Blue = 8'hca;
end 13'h1e8:    begin Red = 8'hfb;    Green = 8'hec;    Blue = 8'hca;
end 13'h1e9:    begin Red = 8'hff;    Green = 8'hea;    Blue = 8'hc8;
end 13'h1ea:    begin Red = 8'he3;    Green = 8'hcc;    Blue = 8'hab;
end 13'h1eb:    begin Red = 8'hfb;    Green = 8'he5;    Blue = 8'hc2;
end 13'h1ec:    begin Red = 8'h9e;    Green = 8'h8a;    Blue = 8'h71;
end 13'h1ed:    begin Red = 8'ha9;    Green = 8'h94;    Blue = 8'h7f;
end 13'h1ee:    begin Red = 8'h84;    Green = 8'h74;    Blue = 8'h5d;
end 13'h1ef:    begin Red = 8'h83;    Green = 8'h70;    Blue = 8'h5b;
end 13'h1f0:    begin Red = 8'hc7;    Green = 8'hb6;    Blue = 8'h97;
end 13'h1f1:    begin Red = 8'hc9;    Green = 8'hb4;    Blue = 8'h98;
end 13'h1f2:    begin Red = 8'ha2;    Green = 8'h8d;    Blue = 8'h79;
end 13'h1f3:    begin Red = 8'h9c;    Green = 8'h89;    Blue = 8'h76;
end 13'h1f4:    begin Red = 8'hde;    Green = 8'hcc;    Blue = 8'hac;
end 13'h1f5:    begin Red = 8'hb8;    Green = 8'ha3;    Blue = 8'h86;
end 13'h1f6:    begin Red = 8'h9b;    Green = 8'h89;    Blue = 8'h6c;
end 13'h1f7:    begin Red = 8'hf9;    Green = 8'he5;    Blue = 8'hbf;
end 13'h1f8:    begin Red = 8'hee;    Green = 8'hdd;    Blue = 8'hb7;
end 13'h1f9:    begin Red = 8'h86;    Green = 8'had;    Blue = 8'h94;
end 13'h1fa:    begin Red = 8'h9c;    Green = 8'haf;    Blue = 8'h96;
end 13'h1fb:    begin Red = 8'h8c;    Green = 8'ha6;    Blue = 8'h82;
end 13'h1fc:    begin Red = 8'hea;    Green = 8'hea;    Blue = 8'heb;
end 13'h1fd:    begin Red = 8'he5;    Green = 8'hea;    Blue = 8'he5;
end 13'h1fe:    begin Red = 8'hed;    Green = 8'hea;    Blue = 8'hef;
end 13'h1ff:    begin Red = 8'hf9;    Green = 8'hfc;    Blue = 8'hfb;
end 13'h200:    begin Red = 8'he4;    Green = 8'heb;    Blue = 8'he9;
end 13'h201:    begin Red = 8'heb;    Green = 8'hf0;    Blue = 8'he8;
end 13'h202:    begin Red = 8'h98;    Green = 8'hb3;    Blue = 8'h92;
end 13'h203:    begin Red = 8'h90;    Green = 8'had;    Blue = 8'h8c;
end 13'h204:    begin Red = 8'h82;    Green = 8'h8c;    Blue = 8'h7e;
end 13'h205:    begin Red = 8'h8d;    Green = 8'hac;    Blue = 8'h87;
end 13'h206:    begin Red = 8'h7e;    Green = 8'h8c;    Blue = 8'h7b;
end 13'h207:    begin Red = 8'h75;    Green = 8'h8d;    Blue = 8'h71;
end 13'h208:    begin Red = 8'h6b;    Green = 8'h82;    Blue = 8'h69;
end 13'h209:    begin Red = 8'h69;    Green = 8'h80;    Blue = 8'h68;
end 13'h20a:    begin Red = 8'h7f;    Green = 8'h94;    Blue = 8'h78;
end 13'h20b:    begin Red = 8'h7a;    Green = 8'h84;    Blue = 8'h76;
end 13'h20c:    begin Red = 8'h6f;    Green = 8'h84;    Blue = 8'h6c;
end 13'h20d:    begin Red = 8'h75;    Green = 8'h88;    Blue = 8'h73;
end 13'h20e:    begin Red = 8'h87;    Green = 8'h9a;    Blue = 8'h87;
end 13'h20f:    begin Red = 8'h6b;    Green = 8'h87;    Blue = 8'h77;
end 13'h210:    begin Red = 8'h70;    Green = 8'h88;    Blue = 8'h6c;
end 13'h211:    begin Red = 8'h6e;    Green = 8'h83;    Blue = 8'h6f;
end 13'h212:    begin Red = 8'h61;    Green = 8'h72;    Blue = 8'h83;
end 13'h213:    begin Red = 8'h46;    Green = 8'h65;    Blue = 8'h69;
end 13'h214:    begin Red = 8'h48;    Green = 8'h66;    Blue = 8'h6d;
end 13'h215:    begin Red = 8'h49;    Green = 8'h61;    Blue = 8'h72;
end 13'h216:    begin Red = 8'h51;    Green = 8'h6c;    Blue = 8'h6e;
end 13'h217:    begin Red = 8'ha8;    Green = 8'ha7;    Blue = 8'h98;
end 13'h218:    begin Red = 8'h71;    Green = 8'h7d;    Blue = 8'h4e;
end 13'h219:    begin Red = 8'h6e;    Green = 8'h78;    Blue = 8'h4c;
end 13'h21a:    begin Red = 8'h6a;    Green = 8'h79;    Blue = 8'h7e;
end 13'h21b:    begin Red = 8'h76;    Green = 8'h7d;    Blue = 8'h4e;
end 13'h21c:    begin Red = 8'h73;    Green = 8'h7f;    Blue = 8'h4b;
end 13'h21d:    begin Red = 8'h88;    Green = 8'h90;    Blue = 8'h5e;
end 13'h21e:    begin Red = 8'h86;    Green = 8'h98;    Blue = 8'h5d;
end 13'h21f:    begin Red = 8'ha1;    Green = 8'hb1;    Blue = 8'h51;
end 13'h220:    begin Red = 8'h66;    Green = 8'h7f;    Blue = 8'h8f;
end 13'h221:    begin Red = 8'h5e;    Green = 8'h7a;    Blue = 8'h7f;
end 13'h222:    begin Red = 8'hf6;    Green = 8'he8;    Blue = 8'hc2;
end 13'h223:    begin Red = 8'h91;    Green = 8'h7f;    Blue = 8'h64;
end 13'h224:    begin Red = 8'hca;    Green = 8'hb8;    Blue = 8'h97;
end 13'h225:    begin Red = 8'hcd;    Green = 8'hb5;    Blue = 8'h98;
end 13'h226:    begin Red = 8'h89;    Green = 8'h7a;    Blue = 8'h60;
end 13'h227:    begin Red = 8'h7d;    Green = 8'h6e;    Blue = 8'h56;
end 13'h228:    begin Red = 8'h8c;    Green = 8'h78;    Blue = 8'h64;
end 13'h229:    begin Red = 8'hb7;    Green = 8'ha6;    Blue = 8'h85;
end 13'h22a:    begin Red = 8'hd2;    Green = 8'hbb;    Blue = 8'ha0;
end 13'h22b:    begin Red = 8'ha3;    Green = 8'h94;    Blue = 8'h78;
end 13'h22c:    begin Red = 8'hc2;    Green = 8'haf;    Blue = 8'h92;
end 13'h22d:    begin Red = 8'h80;    Green = 8'ha9;    Blue = 8'h90;
end 13'h22e:    begin Red = 8'ha0;    Green = 8'hbd;    Blue = 8'h9f;
end 13'h22f:    begin Red = 8'hde;    Green = 8'hdd;    Blue = 8'hd9;
end 13'h230:    begin Red = 8'hd9;    Green = 8'hd8;    Blue = 8'hd6;
end 13'h231:    begin Red = 8'hf9;    Green = 8'hec;    Blue = 8'hf5;
end 13'h232:    begin Red = 8'h89;    Green = 8'h94;    Blue = 8'h86;
end 13'h233:    begin Red = 8'hdb;    Green = 8'hda;    Blue = 8'hd7;
end 13'h234:    begin Red = 8'hd7;    Green = 8'hd6;    Blue = 8'hd5;
end 13'h235:    begin Red = 8'hdf;    Green = 8'hde;    Blue = 8'hdd;
end 13'h236:    begin Red = 8'hdb;    Green = 8'he0;    Blue = 8'hd5;
end 13'h237:    begin Red = 8'h69;    Green = 8'h7d;    Blue = 8'h7d;
end 13'h238:    begin Red = 8'he1;    Green = 8'he2;    Blue = 8'hd8;
end 13'h239:    begin Red = 8'hd2;    Green = 8'hd7;    Blue = 8'hcf;
end 13'h23a:    begin Red = 8'hde;    Green = 8'hdb;    Blue = 8'he2;
end 13'h23b:    begin Red = 8'hf6;    Green = 8'hf9;    Blue = 8'hf3;
end 13'h23c:    begin Red = 8'h4f;    Green = 8'h6c;    Blue = 8'h71;
end 13'h23d:    begin Red = 8'h66;    Green = 8'h81;    Blue = 8'h83;
end 13'h23e:    begin Red = 8'hdd;    Green = 8'hd9;    Blue = 8'hb7;
end 13'h23f:    begin Red = 8'hce;    Green = 8'hce;    Blue = 8'hb1;
end 13'h240:    begin Red = 8'hc2;    Green = 8'hc2;    Blue = 8'hba;
end 13'h241:    begin Red = 8'hb2;    Green = 8'hb2;    Blue = 8'haa;
end 13'h242:    begin Red = 8'h84;    Green = 8'h91;    Blue = 8'h5f;
end 13'h243:    begin Red = 8'h89;    Green = 8'h97;    Blue = 8'h57;
end 13'h244:    begin Red = 8'h69;    Green = 8'h75;    Blue = 8'h48;
end 13'h245:    begin Red = 8'h6d;    Green = 8'h7c;    Blue = 8'h4e;
end 13'h246:    begin Red = 8'h63;    Green = 8'h78;    Blue = 8'h8e;
end 13'h247:    begin Red = 8'h75;    Green = 8'h7e;    Blue = 8'h48;
end 13'h248:    begin Red = 8'h8a;    Green = 8'h98;    Blue = 8'h5f;
end 13'h249:    begin Red = 8'h87;    Green = 8'h94;    Blue = 8'h58;
end 13'h24a:    begin Red = 8'h98;    Green = 8'ha9;    Blue = 8'h59;
end 13'h24b:    begin Red = 8'h67;    Green = 8'h75;    Blue = 8'h83;
end 13'h24c:    begin Red = 8'hd4;    Green = 8'hc5;    Blue = 8'hab;
end 13'h24d:    begin Red = 8'hc0;    Green = 8'had;    Blue = 8'h90;
end 13'h24e:    begin Red = 8'h9f;    Green = 8'h8c;    Blue = 8'h74;
end 13'h24f:    begin Red = 8'ha8;    Green = 8'h93;    Blue = 8'h7c;
end 13'h250:    begin Red = 8'h88;    Green = 8'h78;    Blue = 8'h63;
end 13'h251:    begin Red = 8'hb7;    Green = 8'ha3;    Blue = 8'h8a;
end 13'h252:    begin Red = 8'h95;    Green = 8'h83;    Blue = 8'h69;
end 13'h253:    begin Red = 8'he3;    Green = 8'he2;    Blue = 8'he2;
end 13'h254:    begin Red = 8'he3;    Green = 8'he4;    Blue = 8'hdf;
end 13'h255:    begin Red = 8'he5;    Green = 8'he2;    Blue = 8'hde;
end 13'h256:    begin Red = 8'ha0;    Green = 8'hba;    Blue = 8'h9c;
end 13'h257:    begin Red = 8'h9f;    Green = 8'hba;    Blue = 8'ha0;
end 13'h258:    begin Red = 8'hd2;    Green = 8'hd3;    Blue = 8'hd2;
end 13'h259:    begin Red = 8'hd6;    Green = 8'hdc;    Blue = 8'hd6;
end 13'h25a:    begin Red = 8'hda;    Green = 8'hdb;    Blue = 8'hdd;
end 13'h25b:    begin Red = 8'hf1;    Green = 8'hf2;    Blue = 8'hf6;
end 13'h25c:    begin Red = 8'h6c;    Green = 8'h80;    Blue = 8'h66;
end 13'h25d:    begin Red = 8'h85;    Green = 8'h93;    Blue = 8'h8b;
end 13'h25e:    begin Red = 8'hd9;    Green = 8'hd6;    Blue = 8'hd1;
end 13'h25f:    begin Red = 8'hd6;    Green = 8'hdb;    Blue = 8'hd2;
end 13'h260:    begin Red = 8'hd8;    Green = 8'hdd;    Blue = 8'hd9;
end 13'h261:    begin Red = 8'h3d;    Green = 8'h4e;    Blue = 8'h59;
end 13'h262:    begin Red = 8'h5d;    Green = 8'h69;    Blue = 8'h71;
end 13'h263:    begin Red = 8'hdb;    Green = 8'hd7;    Blue = 8'hb6;
end 13'h264:    begin Red = 8'ha1;    Green = 8'ha0;    Blue = 8'h90;
end 13'h265:    begin Red = 8'ha2;    Green = 8'ha2;    Blue = 8'h8d;
end 13'h266:    begin Red = 8'h8a;    Green = 8'h98;    Blue = 8'h5a;
end 13'h267:    begin Red = 8'h6f;    Green = 8'h73;    Blue = 8'h45;
end 13'h268:    begin Red = 8'h71;    Green = 8'h78;    Blue = 8'h51;
end 13'h269:    begin Red = 8'h73;    Green = 8'h7d;    Blue = 8'h51;
end 13'h26a:    begin Red = 8'h56;    Green = 8'h71;    Blue = 8'h89;
end 13'h26b:    begin Red = 8'hd0;    Green = 8'hc2;    Blue = 8'haf;
end 13'h26c:    begin Red = 8'hff;    Green = 8'hed;    Blue = 8'hca;
end 13'h26d:    begin Red = 8'h88;    Green = 8'h7b;    Blue = 8'h65;
end 13'h26e:    begin Red = 8'ha8;    Green = 8'h97;    Blue = 8'h78;
end 13'h26f:    begin Red = 8'hf9;    Green = 8'hf1;    Blue = 8'hfa;
end 13'h270:    begin Red = 8'he3;    Green = 8'he7;    Blue = 8'hea;
end 13'h271:    begin Red = 8'hd4;    Green = 8'hd4;    Blue = 8'hd4;
end 13'h272:    begin Red = 8'hdb;    Green = 8'hdf;    Blue = 8'hdc;
end 13'h273:    begin Red = 8'hf3;    Green = 8'he7;    Blue = 8'heb;
end 13'h274:    begin Red = 8'hd8;    Green = 8'hd7;    Blue = 8'hdb;
end 13'h275:    begin Red = 8'hf5;    Green = 8'hea;    Blue = 8'hf9;
end 13'h276:    begin Red = 8'h81;    Green = 8'h91;    Blue = 8'h88;
end 13'h277:    begin Red = 8'hd9;    Green = 8'hdb;    Blue = 8'hd0;
end 13'h278:    begin Red = 8'he0;    Green = 8'hd8;    Blue = 8'hd7;
end 13'h279:    begin Red = 8'h3a;    Green = 8'h51;    Blue = 8'h5a;
end 13'h27a:    begin Red = 8'h97;    Green = 8'h95;    Blue = 8'h89;
end 13'h27b:    begin Red = 8'h58;    Green = 8'h67;    Blue = 8'h3b;
end 13'h27c:    begin Red = 8'h5b;    Green = 8'h5d;    Blue = 8'h3e;
end 13'h27d:    begin Red = 8'h5d;    Green = 8'h63;    Blue = 8'h49;
end 13'h27e:    begin Red = 8'h55;    Green = 8'h5c;    Blue = 8'h49;
end 13'h27f:    begin Red = 8'h6f;    Green = 8'h7b;    Blue = 8'h44;
end 13'h280:    begin Red = 8'h9e;    Green = 8'hb1;    Blue = 8'h63;
end 13'h281:    begin Red = 8'h69;    Green = 8'h6c;    Blue = 8'h5f;
end 13'h282:    begin Red = 8'h81;    Green = 8'h8e;    Blue = 8'h55;
end 13'h283:    begin Red = 8'ha0;    Green = 8'hb5;    Blue = 8'h49;
end 13'h284:    begin Red = 8'h9c;    Green = 8'hb0;    Blue = 8'h4a;
end 13'h285:    begin Red = 8'hf1;    Green = 8'hda;    Blue = 8'hbb;
end 13'h286:    begin Red = 8'hce;    Green = 8'hb7;    Blue = 8'h9a;
end 13'h287:    begin Red = 8'h7f;    Green = 8'h6e;    Blue = 8'h5f;
end 13'h288:    begin Red = 8'hba;    Green = 8'hab;    Blue = 8'h8b;
end 13'h289:    begin Red = 8'hf8;    Green = 8'hef;    Blue = 8'hf4;
end 13'h28a:    begin Red = 8'he5;    Green = 8'he5;    Blue = 8'he5;
end 13'h28b:    begin Red = 8'h7f;    Green = 8'h8e;    Blue = 8'h7d;
end 13'h28c:    begin Red = 8'h9b;    Green = 8'hb9;    Blue = 8'h98;
end 13'h28d:    begin Red = 8'he2;    Green = 8'hdf;    Blue = 8'hde;
end 13'h28e:    begin Red = 8'hef;    Green = 8'hed;    Blue = 8'hf2;
end 13'h28f:    begin Red = 8'he9;    Green = 8'hde;    Blue = 8'hd9;
end 13'h290:    begin Red = 8'h6a;    Green = 8'h84;    Blue = 8'h6d;
end 13'h291:    begin Red = 8'hdf;    Green = 8'he3;    Blue = 8'he0;
end 13'h292:    begin Red = 8'hcf;    Green = 8'hcf;    Blue = 8'hc9;
end 13'h293:    begin Red = 8'hef;    Green = 8'he6;    Blue = 8'heb;
end 13'h294:    begin Red = 8'hd8;    Green = 8'hd6;    Blue = 8'hcd;
end 13'h295:    begin Red = 8'h72;    Green = 8'h81;    Blue = 8'h70;
end 13'h296:    begin Red = 8'h6e;    Green = 8'h7c;    Blue = 8'h6c;
end 13'h297:    begin Red = 8'hd6;    Green = 8'hd5;    Blue = 8'hd2;
end 13'h298:    begin Red = 8'hf2;    Green = 8'heb;    Blue = 8'hef;
end 13'h299:    begin Red = 8'h75;    Green = 8'h7e;    Blue = 8'h73;
end 13'h29a:    begin Red = 8'hd7;    Green = 8'hd3;    Blue = 8'hb5;
end 13'h29b:    begin Red = 8'hcc;    Green = 8'hcc;    Blue = 8'haf;
end 13'h29c:    begin Red = 8'h55;    Green = 8'h5d;    Blue = 8'h40;
end 13'h29d:    begin Red = 8'h72;    Green = 8'h7c;    Blue = 8'h54;
end 13'h29e:    begin Red = 8'h70;    Green = 8'h7a;    Blue = 8'h4f;
end 13'h29f:    begin Red = 8'h6f;    Green = 8'h7e;    Blue = 8'h51;
end 13'h2a0:    begin Red = 8'h5e;    Green = 8'h61;    Blue = 8'h3b;
end 13'h2a1:    begin Red = 8'h55;    Green = 8'h67;    Blue = 8'h40;
end 13'h2a2:    begin Red = 8'h58;    Green = 8'h60;    Blue = 8'h42;
end 13'h2a3:    begin Red = 8'h7b;    Green = 8'h88;    Blue = 8'h4f;
end 13'h2a4:    begin Red = 8'h78;    Green = 8'h84;    Blue = 8'h50;
end 13'h2a5:    begin Red = 8'h67;    Green = 8'h5d;    Blue = 8'h61;
end 13'h2a6:    begin Red = 8'h6c;    Green = 8'h6a;    Blue = 8'h66;
end 13'h2a7:    begin Red = 8'h80;    Green = 8'h8d;    Blue = 8'h5c;
end 13'h2a8:    begin Red = 8'ha8;    Green = 8'hbc;    Blue = 8'h3b;
end 13'h2a9:    begin Red = 8'ha8;    Green = 8'hbb;    Blue = 8'h34;
end 13'h2aa:    begin Red = 8'hba;    Green = 8'hd2;    Blue = 8'h3a;
end 13'h2ab:    begin Red = 8'hca;    Green = 8'hde;    Blue = 8'h34;
end 13'h2ac:    begin Red = 8'hef;    Green = 8'hd9;    Blue = 8'hb7;
end 13'h2ad:    begin Red = 8'h97;    Green = 8'h85;    Blue = 8'h65;
end 13'h2ae:    begin Red = 8'hac;    Green = 8'h99;    Blue = 8'h7b;
end 13'h2af:    begin Red = 8'h81;    Green = 8'h6f;    Blue = 8'h62;
end 13'h2b0:    begin Red = 8'h84;    Green = 8'h70;    Blue = 8'h60;
end 13'h2b1:    begin Red = 8'h77;    Green = 8'h64;    Blue = 8'h4f;
end 13'h2b2:    begin Red = 8'hb9;    Green = 8'ha5;    Blue = 8'h8d;
end 13'h2b3:    begin Red = 8'hbd;    Green = 8'hac;    Blue = 8'h8c;
end 13'h2b4:    begin Red = 8'h7d;    Green = 8'h6b;    Blue = 8'h5e;
end 13'h2b5:    begin Red = 8'h7e;    Green = 8'h6c;    Blue = 8'h5a;
end 13'h2b6:    begin Red = 8'h7b;    Green = 8'h6d;    Blue = 8'h59;
end 13'h2b7:    begin Red = 8'ha7;    Green = 8'h92;    Blue = 8'h81;
end 13'h2b8:    begin Red = 8'hbb;    Green = 8'ha4;    Blue = 8'h84;
end 13'h2b9:    begin Red = 8'hf6;    Green = 8'hdc;    Blue = 8'hc0;
end 13'h2ba:    begin Red = 8'he1;    Green = 8'he6;    Blue = 8'he1;
end 13'h2bb:    begin Red = 8'hf6;    Green = 8'hee;    Blue = 8'hf2;
end 13'h2bc:    begin Red = 8'hf6;    Green = 8'hf2;    Blue = 8'hf1;
end 13'h2bd:    begin Red = 8'he2;    Green = 8'he0;    Blue = 8'hda;
end 13'h2be:    begin Red = 8'h9d;    Green = 8'hb7;    Blue = 8'ha4;
end 13'h2bf:    begin Red = 8'h95;    Green = 8'hb5;    Blue = 8'h99;
end 13'h2c0:    begin Red = 8'h88;    Green = 8'ha9;    Blue = 8'h8e;
end 13'h2c1:    begin Red = 8'h80;    Green = 8'ha7;    Blue = 8'h7f;
end 13'h2c2:    begin Red = 8'hf0;    Green = 8'hec;    Blue = 8'he7;
end 13'h2c3:    begin Red = 8'hee;    Green = 8'hf1;    Blue = 8'hea;
end 13'h2c4:    begin Red = 8'ha5;    Green = 8'hb9;    Blue = 8'ha1;
end 13'h2c5:    begin Red = 8'h78;    Green = 8'h83;    Blue = 8'h71;
end 13'h2c6:    begin Red = 8'hfd;    Green = 8'heb;    Blue = 8'hf5;
end 13'h2c7:    begin Red = 8'hf4;    Green = 8'hf0;    Blue = 8'hf6;
end 13'h2c8:    begin Red = 8'hd6;    Green = 8'hd2;    Blue = 8'hd0;
end 13'h2c9:    begin Red = 8'hce;    Green = 8'hd3;    Blue = 8'hca;
end 13'h2ca:    begin Red = 8'hd5;    Green = 8'hd1;    Blue = 8'hcc;
end 13'h2cb:    begin Red = 8'h6f;    Green = 8'h81;    Blue = 8'h75;
end 13'h2cc:    begin Red = 8'hce;    Green = 8'hd7;    Blue = 8'hcc;
end 13'h2cd:    begin Red = 8'h70;    Green = 8'h7f;    Blue = 8'h6d;
end 13'h2ce:    begin Red = 8'h6d;    Green = 8'h87;    Blue = 8'h68;
end 13'h2cf:    begin Red = 8'h62;    Green = 8'h7d;    Blue = 8'h67;
end 13'h2d0:    begin Red = 8'hd6;    Green = 8'hce;    Blue = 8'hcf;
end 13'h2d1:    begin Red = 8'h5c;    Green = 8'h67;    Blue = 8'h6e;
end 13'h2d2:    begin Red = 8'h9d;    Green = 8'h9c;    Blue = 8'h8e;
end 13'h2d3:    begin Red = 8'h78;    Green = 8'h81;    Blue = 8'h4d;
end 13'h2d4:    begin Red = 8'h5d;    Green = 8'h64;    Blue = 8'h43;
end 13'h2d5:    begin Red = 8'h78;    Green = 8'h7d;    Blue = 8'h52;
end 13'h2d6:    begin Red = 8'h6b;    Green = 8'h69;    Blue = 8'h5b;
end 13'h2d7:    begin Red = 8'h70;    Green = 8'h70;    Blue = 8'h53;
end 13'h2d8:    begin Red = 8'h90;    Green = 8'h9b;    Blue = 8'h56;
end 13'h2d9:    begin Red = 8'h89;    Green = 8'h96;    Blue = 8'h62;
end 13'h2da:    begin Red = 8'ha3;    Green = 8'hb7;    Blue = 8'h41;
end 13'h2db:    begin Red = 8'h98;    Green = 8'hab;    Blue = 8'h43;
end 13'h2dc:    begin Red = 8'haa;    Green = 8'hc0;    Blue = 8'h4d;
end 13'h2dd:    begin Red = 8'hc2;    Green = 8'hce;    Blue = 8'h3c;
end 13'h2de:    begin Red = 8'h94;    Green = 8'h82;    Blue = 8'h63;
end 13'h2df:    begin Red = 8'hb5;    Green = 8'ha2;    Blue = 8'h87;
end 13'h2e0:    begin Red = 8'h88;    Green = 8'h77;    Blue = 8'h5e;
end 13'h2e1:    begin Red = 8'hc0;    Green = 8'haa;    Blue = 8'h8b;
end 13'h2e2:    begin Red = 8'hd3;    Green = 8'hb9;    Blue = 8'h9d;
end 13'h2e3:    begin Red = 8'hf6;    Green = 8'hed;    Blue = 8'hf8;
end 13'h2e4:    begin Red = 8'he8;    Green = 8'hdf;    Blue = 8'he2;
end 13'h2e5:    begin Red = 8'h6a;    Green = 8'h7c;    Blue = 8'h69;
end 13'h2e6:    begin Red = 8'h72;    Green = 8'h89;    Blue = 8'h71;
end 13'h2e7:    begin Red = 8'h61;    Green = 8'h7a;    Blue = 8'h75;
end 13'h2e8:    begin Red = 8'hd5;    Green = 8'hd1;    Blue = 8'hb3;
end 13'h2e9:    begin Red = 8'hca;    Green = 8'hc8;    Blue = 8'haf;
end 13'h2ea:    begin Red = 8'hbc;    Green = 8'hbc;    Blue = 8'hb4;
end 13'h2eb:    begin Red = 8'h8b;    Green = 8'h8c;    Blue = 8'h79;
end 13'h2ec:    begin Red = 8'ha2;    Green = 8'ha4;    Blue = 8'h9d;
end 13'h2ed:    begin Red = 8'hb1;    Green = 8'hb3;    Blue = 8'ha4;
end 13'h2ee:    begin Red = 8'had;    Green = 8'hb0;    Blue = 8'h9e;
end 13'h2ef:    begin Red = 8'h5c;    Green = 8'h63;    Blue = 8'h3e;
end 13'h2f0:    begin Red = 8'h5a;    Green = 8'h63;    Blue = 8'h3b;
end 13'h2f1:    begin Red = 8'h71;    Green = 8'h71;    Blue = 8'h61;
end 13'h2f2:    begin Red = 8'h71;    Green = 8'h71;    Blue = 8'h58;
end 13'h2f3:    begin Red = 8'h6c;    Green = 8'h6f;    Blue = 8'h5a;
end 13'h2f4:    begin Red = 8'h81;    Green = 8'h93;    Blue = 8'h57;
end 13'h2f5:    begin Red = 8'h88;    Green = 8'h96;    Blue = 8'h4b;
end 13'h2f6:    begin Red = 8'h66;    Green = 8'h80;    Blue = 8'h7c;
end 13'h2f7:    begin Red = 8'h5f;    Green = 8'h79;    Blue = 8'h85;
end 13'h2f8:    begin Red = 8'h89;    Green = 8'h78;    Blue = 8'h68;
end 13'h2f9:    begin Red = 8'hb9;    Green = 8'ha6;    Blue = 8'h89;
end 13'h2fa:    begin Red = 8'h96;    Green = 8'hac;    Blue = 8'h5a;
end 13'h2fb:    begin Red = 8'h98;    Green = 8'hbc;    Blue = 8'ha3;
end 13'h2fc:    begin Red = 8'hf4;    Green = 8'hec;    Blue = 8'hf5;
end 13'h2fd:    begin Red = 8'hda;    Green = 8'he3;    Blue = 8'he0;
end 13'h2fe:    begin Red = 8'h81;    Green = 8'h96;    Blue = 8'h82;
end 13'h2ff:    begin Red = 8'h6f;    Green = 8'h89;    Blue = 8'h74;
end 13'h300:    begin Red = 8'hf0;    Green = 8'hed;    Blue = 8'hec;
end 13'h301:    begin Red = 8'hd1;    Green = 8'hce;    Blue = 8'hcb;
end 13'h302:    begin Red = 8'hce;    Green = 8'hce;    Blue = 8'hc6;
end 13'h303:    begin Red = 8'h92;    Green = 8'h91;    Blue = 8'h83;
end 13'h304:    begin Red = 8'h8e;    Green = 8'h8c;    Blue = 8'h80;
end 13'h305:    begin Red = 8'h94;    Green = 8'ha3;    Blue = 8'h5a;
end 13'h306:    begin Red = 8'haf;    Green = 8'hb0;    Blue = 8'hb3;
end 13'h307:    begin Red = 8'h52;    Green = 8'h5a;    Blue = 8'h3f;
end 13'h308:    begin Red = 8'h78;    Green = 8'h7e;    Blue = 8'h5d;
end 13'h309:    begin Red = 8'h77;    Green = 8'h7d;    Blue = 8'h56;
end 13'h30a:    begin Red = 8'h59;    Green = 8'h5e;    Blue = 8'h44;
end 13'h30b:    begin Red = 8'h59;    Green = 8'h5f;    Blue = 8'h36;
end 13'h30c:    begin Red = 8'h67;    Green = 8'h65;    Blue = 8'h5d;
end 13'h30d:    begin Red = 8'h68;    Green = 8'h62;    Blue = 8'h5c;
end 13'h30e:    begin Red = 8'h69;    Green = 8'h65;    Blue = 8'h61;
end 13'h30f:    begin Red = 8'h80;    Green = 8'h98;    Blue = 8'h58;
end 13'h310:    begin Red = 8'h8e;    Green = 8'h91;    Blue = 8'h54;
end 13'h311:    begin Red = 8'h8b;    Green = 8'ha0;    Blue = 8'h56;
end 13'h312:    begin Red = 8'h5b;    Green = 8'h77;    Blue = 8'h88;
end 13'h313:    begin Red = 8'h65;    Green = 8'h78;    Blue = 8'h80;
end 13'h314:    begin Red = 8'h6c;    Green = 8'h7b;    Blue = 8'h83;
end 13'h315:    begin Red = 8'hc8;    Green = 8'hb0;    Blue = 8'h9b;
end 13'h316:    begin Red = 8'hc6;    Green = 8'hb1;    Blue = 8'h95;
end 13'h317:    begin Red = 8'hc5;    Green = 8'hb3;    Blue = 8'h9a;
end 13'h318:    begin Red = 8'hd0;    Green = 8'hab;    Blue = 8'h9b;
end 13'h319:    begin Red = 8'h8d;    Green = 8'h75;    Blue = 8'h66;
end 13'h31a:    begin Red = 8'h89;    Green = 8'h71;    Blue = 8'h62;
end 13'h31b:    begin Red = 8'hb2;    Green = 8'h99;    Blue = 8'h88;
end 13'h31c:    begin Red = 8'hc1;    Green = 8'ha5;    Blue = 8'h96;
end 13'h31d:    begin Red = 8'hc6;    Green = 8'ha5;    Blue = 8'h8d;
end 13'h31e:    begin Red = 8'hd6;    Green = 8'hb7;    Blue = 8'ha7;
end 13'h31f:    begin Red = 8'h92;    Green = 8'h87;    Blue = 8'h68;
end 13'h320:    begin Red = 8'hed;    Green = 8'he1;    Blue = 8'hba;
end 13'h321:    begin Red = 8'had;    Green = 8'h92;    Blue = 8'h7d;
end 13'h322:    begin Red = 8'hfe;    Green = 8'heb;    Blue = 8'hd5;
end 13'h323:    begin Red = 8'hff;    Green = 8'hee;    Blue = 8'hd8;
end 13'h324:    begin Red = 8'h90;    Green = 8'ha8;    Blue = 8'h61;
end 13'h325:    begin Red = 8'h9b;    Green = 8'ha8;    Blue = 8'h54;
end 13'h326:    begin Red = 8'ha0;    Green = 8'hb7;    Blue = 8'ha8;
end 13'h327:    begin Red = 8'hf2;    Green = 8'hea;    Blue = 8'hf3;
end 13'h328:    begin Red = 8'he1;    Green = 8'hd9;    Blue = 8'hde;
end 13'h329:    begin Red = 8'he2;    Green = 8'hdb;    Blue = 8'hdc;
end 13'h32a:    begin Red = 8'h8c;    Green = 8'hab;    Blue = 8'h8a;
end 13'h32b:    begin Red = 8'h70;    Green = 8'h8a;    Blue = 8'h68;
end 13'h32c:    begin Red = 8'he4;    Green = 8'hdd;    Blue = 8'he1;
end 13'h32d:    begin Red = 8'hd4;    Green = 8'hd9;    Blue = 8'hd9;
end 13'h32e:    begin Red = 8'h72;    Green = 8'h81;    Blue = 8'h6b;
end 13'h32f:    begin Red = 8'h60;    Green = 8'h71;    Blue = 8'h8f;
end 13'h330:    begin Red = 8'h5e;    Green = 8'h73;    Blue = 8'h80;
end 13'h331:    begin Red = 8'h9c;    Green = 8'h9f;    Blue = 8'h89;
end 13'h332:    begin Red = 8'ha0;    Green = 8'h9d;    Blue = 8'h91;
end 13'h333:    begin Red = 8'hbe;    Green = 8'hbb;    Blue = 8'hbb;
end 13'h334:    begin Red = 8'hb5;    Green = 8'hb3;    Blue = 8'hb6;
end 13'h335:    begin Red = 8'hbc;    Green = 8'hc0;    Blue = 8'hb0;
end 13'h336:    begin Red = 8'hc5;    Green = 8'hc3;    Blue = 8'hc7;
end 13'h337:    begin Red = 8'hc3;    Green = 8'hc1;    Blue = 8'hc3;
end 13'h338:    begin Red = 8'hbb;    Green = 8'hbe;    Blue = 8'ha8;
end 13'h339:    begin Red = 8'h9b;    Green = 8'h97;    Blue = 8'h94;
end 13'h33a:    begin Red = 8'h91;    Green = 8'h8e;    Blue = 8'h87;
end 13'h33b:    begin Red = 8'haf;    Green = 8'hac;    Blue = 8'hbf;
end 13'h33c:    begin Red = 8'h5c;    Green = 8'h60;    Blue = 8'h4e;
end 13'h33d:    begin Red = 8'h62;    Green = 8'h69;    Blue = 8'h4a;
end 13'h33e:    begin Red = 8'h83;    Green = 8'h91;    Blue = 8'h56;
end 13'h33f:    begin Red = 8'h81;    Green = 8'h83;    Blue = 8'h63;
end 13'h340:    begin Red = 8'h80;    Green = 8'h80;    Blue = 8'h58;
end 13'h341:    begin Red = 8'h82;    Green = 8'h7f;    Blue = 8'h61;
end 13'h342:    begin Red = 8'h7f;    Green = 8'h7d;    Blue = 8'h59;
end 13'h343:    begin Red = 8'h61;    Green = 8'h7a;    Blue = 8'h70;
end 13'h344:    begin Red = 8'h88;    Green = 8'h76;    Blue = 8'h6b;
end 13'h345:    begin Red = 8'h91;    Green = 8'h78;    Blue = 8'h62;
end 13'h346:    begin Red = 8'haf;    Green = 8'h92;    Blue = 8'h85;
end 13'h347:    begin Red = 8'h68;    Green = 8'h80;    Blue = 8'h4d;
end 13'h348:    begin Red = 8'h65;    Green = 8'h74;    Blue = 8'h42;
end 13'h349:    begin Red = 8'h85;    Green = 8'h96;    Blue = 8'h57;
end 13'h34a:    begin Red = 8'hc8;    Green = 8'hab;    Blue = 8'h9c;
end 13'h34b:    begin Red = 8'hdd;    Green = 8'hbc;    Blue = 8'hab;
end 13'h34c:    begin Red = 8'hed;    Green = 8'hde;    Blue = 8'hb3;
end 13'h34d:    begin Red = 8'h91;    Green = 8'h81;    Blue = 8'h67;
end 13'h34e:    begin Red = 8'hff;    Green = 8'hef;    Blue = 8'hd4;
end 13'h34f:    begin Red = 8'h6c;    Green = 8'h78;    Blue = 8'h46;
end 13'h350:    begin Red = 8'h97;    Green = 8'ha6;    Blue = 8'h51;
end 13'h351:    begin Red = 8'h8f;    Green = 8'hac;    Blue = 8'h57;
end 13'h352:    begin Red = 8'h9b;    Green = 8'hba;    Blue = 8'ha6;
end 13'h353:    begin Red = 8'he1;    Green = 8'hdf;    Blue = 8'he2;
end 13'h354:    begin Red = 8'he1;    Green = 8'he1;    Blue = 8'he7;
end 13'h355:    begin Red = 8'hd5;    Green = 8'hdc;    Blue = 8'hdb;
end 13'h356:    begin Red = 8'hde;    Green = 8'he0;    Blue = 8'hdf;
end 13'h357:    begin Red = 8'hed;    Green = 8'he5;    Blue = 8'he8;
end 13'h358:    begin Red = 8'h86;    Green = 8'h91;    Blue = 8'h7d;
end 13'h359:    begin Red = 8'h66;    Green = 8'h86;    Blue = 8'h69;
end 13'h35a:    begin Red = 8'hce;    Green = 8'hc8;    Blue = 8'hc7;
end 13'h35b:    begin Red = 8'hca;    Green = 8'hc9;    Blue = 8'hc6;
end 13'h35c:    begin Red = 8'hdc;    Green = 8'hd7;    Blue = 8'hd9;
end 13'h35d:    begin Red = 8'hcf;    Green = 8'hd4;    Blue = 8'hd4;
end 13'h35e:    begin Red = 8'hcb;    Green = 8'hca;    Blue = 8'hc9;
end 13'h35f:    begin Red = 8'h6e;    Green = 8'h7f;    Blue = 8'h73;
end 13'h360:    begin Red = 8'h88;    Green = 8'h92;    Blue = 8'h8c;
end 13'h361:    begin Red = 8'hd1;    Green = 8'hcd;    Blue = 8'haf;
end 13'h362:    begin Red = 8'hc3;    Green = 8'hc5;    Blue = 8'ha5;
end 13'h363:    begin Red = 8'h9e;    Green = 8'h9f;    Blue = 8'h85;
end 13'h364:    begin Red = 8'h82;    Green = 8'h95;    Blue = 8'h49;
end 13'h365:    begin Red = 8'h8f;    Green = 8'h92;    Blue = 8'h7e;
end 13'h366:    begin Red = 8'h6c;    Green = 8'h7b;    Blue = 8'h40;
end 13'h367:    begin Red = 8'hc7;    Green = 8'hc1;    Blue = 8'hcb;
end 13'h368:    begin Red = 8'hbb;    Green = 8'hbb;    Blue = 8'had;
end 13'h369:    begin Red = 8'h7a;    Green = 8'h8f;    Blue = 8'h40;
end 13'h36a:    begin Red = 8'hb7;    Green = 8'hbb;    Blue = 8'haf;
end 13'h36b:    begin Red = 8'h87;    Green = 8'h90;    Blue = 8'h51;
end 13'h36c:    begin Red = 8'h95;    Green = 8'had;    Blue = 8'h54;
end 13'h36d:    begin Red = 8'h9a;    Green = 8'hac;    Blue = 8'h65;
end 13'h36e:    begin Red = 8'h88;    Green = 8'h94;    Blue = 8'h5f;
end 13'h36f:    begin Red = 8'h9c;    Green = 8'hac;    Blue = 8'h61;
end 13'h370:    begin Red = 8'hae;    Green = 8'haf;    Blue = 8'haf;
end 13'h371:    begin Red = 8'h86;    Green = 8'h93;    Blue = 8'h61;
end 13'h372:    begin Red = 8'h72;    Green = 8'h72;    Blue = 8'h5c;
end 13'h373:    begin Red = 8'h72;    Green = 8'h6c;    Blue = 8'h63;
end 13'h374:    begin Red = 8'h76;    Green = 8'h71;    Blue = 8'h69;
end 13'h375:    begin Red = 8'h79;    Green = 8'h72;    Blue = 8'h65;
end 13'h376:    begin Red = 8'h77;    Green = 8'h6f;    Blue = 8'h67;
end 13'h377:    begin Red = 8'h8b;    Green = 8'h92;    Blue = 8'h5d;
end 13'h378:    begin Red = 8'h80;    Green = 8'h80;    Blue = 8'h5f;
end 13'h379:    begin Red = 8'h85;    Green = 8'h7c;    Blue = 8'h67;
end 13'h37a:    begin Red = 8'haf;    Green = 8'haf;    Blue = 8'h4e;
end 13'h37b:    begin Red = 8'ha7;    Green = 8'ha9;    Blue = 8'h54;
end 13'h37c:    begin Red = 8'hac;    Green = 8'ha9;    Blue = 8'h55;
end 13'h37d:    begin Red = 8'haf;    Green = 8'ha6;    Blue = 8'h4d;
end 13'h37e:    begin Red = 8'hac;    Green = 8'hac;    Blue = 8'h4d;
end 13'h37f:    begin Red = 8'haa;    Green = 8'hac;    Blue = 8'h3e;
end 13'h380:    begin Red = 8'hc7;    Green = 8'hae;    Blue = 8'h4a;
end 13'h381:    begin Red = 8'h94;    Green = 8'h7f;    Blue = 8'h6b;
end 13'h382:    begin Red = 8'h94;    Green = 8'h7e;    Blue = 8'h67;
end 13'h383:    begin Red = 8'hcb;    Green = 8'hb4;    Blue = 8'h94;
end 13'h384:    begin Red = 8'hca;    Green = 8'hb5;    Blue = 8'h9b;
end 13'h385:    begin Red = 8'haf;    Green = 8'h9b;    Blue = 8'h82;
end 13'h386:    begin Red = 8'h82;    Green = 8'h9b;    Blue = 8'h50;
end 13'h387:    begin Red = 8'h85;    Green = 8'h98;    Blue = 8'h52;
end 13'h388:    begin Red = 8'h64;    Green = 8'h6f;    Blue = 8'h40;
end 13'h389:    begin Red = 8'h65;    Green = 8'h76;    Blue = 8'h3f;
end 13'h38a:    begin Red = 8'h94;    Green = 8'h99;    Blue = 8'h5e;
end 13'h38b:    begin Red = 8'h6b;    Green = 8'h79;    Blue = 8'h4b;
end 13'h38c:    begin Red = 8'h5d;    Green = 8'h73;    Blue = 8'h44;
end 13'h38d:    begin Red = 8'h61;    Green = 8'h70;    Blue = 8'h3d;
end 13'h38e:    begin Red = 8'h7f;    Green = 8'h8c;    Blue = 8'h51;
end 13'h38f:    begin Red = 8'h77;    Green = 8'h89;    Blue = 8'h48;
end 13'h390:    begin Red = 8'h51;    Green = 8'h64;    Blue = 8'h34;
end 13'h391:    begin Red = 8'h68;    Green = 8'h78;    Blue = 8'h3d;
end 13'h392:    begin Red = 8'h5a;    Green = 8'h6b;    Blue = 8'h36;
end 13'h393:    begin Red = 8'h83;    Green = 8'h8e;    Blue = 8'h5d;
end 13'h394:    begin Red = 8'ha4;    Green = 8'hb7;    Blue = 8'h5d;
end 13'h395:    begin Red = 8'h9a;    Green = 8'hbb;    Blue = 8'haa;
end 13'h396:    begin Red = 8'h9c;    Green = 8'hb7;    Blue = 8'hae;
end 13'h397:    begin Red = 8'hef;    Green = 8'he7;    Blue = 8'hf0;
end 13'h398:    begin Red = 8'hd5;    Green = 8'hd5;    Blue = 8'hce;
end 13'h399:    begin Red = 8'hd8;    Green = 8'hde;    Blue = 8'he1;
end 13'h39a:    begin Red = 8'he6;    Green = 8'he4;    Blue = 8'hea;
end 13'h39b:    begin Red = 8'hd5;    Green = 8'hd9;    Blue = 8'hd0;
end 13'h39c:    begin Red = 8'hdb;    Green = 8'hd5;    Blue = 8'hd3;
end 13'h39d:    begin Red = 8'he7;    Green = 8'hdd;    Blue = 8'he4;
end 13'h39e:    begin Red = 8'hcb;    Green = 8'hc5;    Blue = 8'hc3;
end 13'h39f:    begin Red = 8'hd2;    Green = 8'hcd;    Blue = 8'hce;
end 13'h3a0:    begin Red = 8'hcc;    Green = 8'hd1;    Blue = 8'hd1;
end 13'h3a1:    begin Red = 8'hd0;    Green = 8'hd0;    Blue = 8'hd0;
end 13'h3a2:    begin Red = 8'h70;    Green = 8'h80;    Blue = 8'h69;
end 13'h3a3:    begin Red = 8'h85;    Green = 8'h8d;    Blue = 8'h87;
end 13'h3a4:    begin Red = 8'h88;    Green = 8'h9b;    Blue = 8'h80;
end 13'h3a5:    begin Red = 8'hcf;    Green = 8'hcb;    Blue = 8'had;
end 13'h3a6:    begin Red = 8'hc5;    Green = 8'hc5;    Blue = 8'haa;
end 13'h3a7:    begin Red = 8'h9b;    Green = 8'h9b;    Blue = 8'h84;
end 13'h3a8:    begin Red = 8'h83;    Green = 8'h8e;    Blue = 8'h49;
end 13'h3a9:    begin Red = 8'h81;    Green = 8'h91;    Blue = 8'h4e;
end 13'h3aa:    begin Red = 8'h84;    Green = 8'h95;    Blue = 8'h5a;
end 13'h3ab:    begin Red = 8'h67;    Green = 8'h76;    Blue = 8'h43;
end 13'h3ac:    begin Red = 8'h8d;    Green = 8'h9b;    Blue = 8'h5f;
end 13'h3ad:    begin Red = 8'h63;    Green = 8'h6c;    Blue = 8'h36;
end 13'h3ae:    begin Red = 8'h7c;    Green = 8'h90;    Blue = 8'h58;
end 13'h3af:    begin Red = 8'h76;    Green = 8'h90;    Blue = 8'h42;
end 13'h3b0:    begin Red = 8'h75;    Green = 8'h88;    Blue = 8'h35;
end 13'h3b1:    begin Red = 8'hb3;    Green = 8'hb4;    Blue = 8'ha7;
end 13'h3b2:    begin Red = 8'hc6;    Green = 8'hc5;    Blue = 8'hc9;
end 13'h3b3:    begin Red = 8'h61;    Green = 8'h73;    Blue = 8'h39;
end 13'h3b4:    begin Red = 8'h81;    Green = 8'h92;    Blue = 8'h5b;
end 13'h3b5:    begin Red = 8'h9f;    Green = 8'hb3;    Blue = 8'h5c;
end 13'h3b6:    begin Red = 8'h8f;    Green = 8'h82;    Blue = 8'h83;
end 13'h3b7:    begin Red = 8'h81;    Green = 8'h7d;    Blue = 8'h80;
end 13'h3b8:    begin Red = 8'ha7;    Green = 8'ha3;    Blue = 8'ha8;
end 13'h3b9:    begin Red = 8'hac;    Green = 8'hac;    Blue = 8'ha8;
end 13'h3ba:    begin Red = 8'h6f;    Green = 8'h6b;    Blue = 8'h5c;
end 13'h3bb:    begin Red = 8'h67;    Green = 8'h6a;    Blue = 8'h56;
end 13'h3bc:    begin Red = 8'h6d;    Green = 8'h6d;    Blue = 8'h57;
end 13'h3bd:    begin Red = 8'h6a;    Green = 8'h68;    Blue = 8'h64;
end 13'h3be:    begin Red = 8'h60;    Green = 8'h60;    Blue = 8'h60;
end 13'h3bf:    begin Red = 8'h7e;    Green = 8'h88;    Blue = 8'h5d;
end 13'h3c0:    begin Red = 8'h80;    Green = 8'h74;    Blue = 8'h65;
end 13'h3c1:    begin Red = 8'h86;    Green = 8'h7b;    Blue = 8'h5d;
end 13'h3c2:    begin Red = 8'hb3;    Green = 8'hac;    Blue = 8'h4e;
end 13'h3c3:    begin Red = 8'had;    Green = 8'ha7;    Blue = 8'h50;
end 13'h3c4:    begin Red = 8'ha9;    Green = 8'ha1;    Blue = 8'h54;
end 13'h3c5:    begin Red = 8'ha3;    Green = 8'ha2;    Blue = 8'h51;
end 13'h3c6:    begin Red = 8'ha0;    Green = 8'ha4;    Blue = 8'h4e;
end 13'h3c7:    begin Red = 8'hb1;    Green = 8'ha8;    Blue = 8'h44;
end 13'h3c8:    begin Red = 8'h4e;    Green = 8'h6c;    Blue = 8'h94;
end 13'h3c9:    begin Red = 8'h57;    Green = 8'h71;    Blue = 8'h90;
end 13'h3ca:    begin Red = 8'h57;    Green = 8'h74;    Blue = 8'h87;
end 13'h3cb:    begin Red = 8'hf4;    Green = 8'he0;    Blue = 8'hc0;
end 13'h3cc:    begin Red = 8'h90;    Green = 8'h7d;    Blue = 8'h61;
end 13'h3cd:    begin Red = 8'hd4;    Green = 8'hbe;    Blue = 8'h9e;
end 13'h3ce:    begin Red = 8'hc3;    Green = 8'haf;    Blue = 8'h9b;
end 13'h3cf:    begin Red = 8'h74;    Green = 8'h91;    Blue = 8'h51;
end 13'h3d0:    begin Red = 8'h91;    Green = 8'h9e;    Blue = 8'h64;
end 13'h3d1:    begin Red = 8'hff;    Green = 8'hfd;    Blue = 8'hdd;
end 13'h3d2:    begin Red = 8'h5f;    Green = 8'h70;    Blue = 8'h41;
end 13'h3d3:    begin Red = 8'h7b;    Green = 8'h8d;    Blue = 8'h4c;
end 13'h3d4:    begin Red = 8'h6c;    Green = 8'h84;    Blue = 8'h3c;
end 13'h3d5:    begin Red = 8'h84;    Green = 8'h9d;    Blue = 8'h46;
end 13'h3d6:    begin Red = 8'h81;    Green = 8'h98;    Blue = 8'h4e;
end 13'h3d7:    begin Red = 8'h98;    Green = 8'hb7;    Blue = 8'h9e;
end 13'h3d8:    begin Red = 8'hed;    Green = 8'he5;    Blue = 8'hed;
end 13'h3d9:    begin Red = 8'h91;    Green = 8'haf;    Blue = 8'h90;
end 13'h3da:    begin Red = 8'hd9;    Green = 8'hd3;    Blue = 8'hce;
end 13'h3db:    begin Red = 8'h6a;    Green = 8'h8b;    Blue = 8'h6b;
end 13'h3dc:    begin Red = 8'h62;    Green = 8'h7f;    Blue = 8'h61;
end 13'h3dd:    begin Red = 8'h8d;    Green = 8'hae;    Blue = 8'h8b;
end 13'h3de:    begin Red = 8'he0;    Green = 8'hd2;    Blue = 8'hd9;
end 13'h3df:    begin Red = 8'hed;    Green = 8'he8;    Blue = 8'he3;
end 13'h3e0:    begin Red = 8'h7d;    Green = 8'h8c;    Blue = 8'h77;
end 13'h3e1:    begin Red = 8'hc6;    Green = 8'hc5;    Blue = 8'hc1;
end 13'h3e2:    begin Red = 8'h8a;    Green = 8'h9a;    Blue = 8'h84;
end 13'h3e3:    begin Red = 8'h71;    Green = 8'h8e;    Blue = 8'h6b;
end 13'h3e4:    begin Red = 8'h62;    Green = 8'h80;    Blue = 8'h65;
end 13'h3e5:    begin Red = 8'h55;    Green = 8'h6f;    Blue = 8'h7b;
end 13'h3e6:    begin Red = 8'hc7;    Green = 8'hc5;    Blue = 8'ha6;
end 13'h3e7:    begin Red = 8'h82;    Green = 8'h92;    Blue = 8'h4b;
end 13'h3e8:    begin Red = 8'h83;    Green = 8'h95;    Blue = 8'h4e;
end 13'h3e9:    begin Red = 8'h90;    Green = 8'h9e;    Blue = 8'h5a;
end 13'h3ea:    begin Red = 8'h69;    Green = 8'h74;    Blue = 8'h4d;
end 13'h3eb:    begin Red = 8'h69;    Green = 8'h75;    Blue = 8'h3f;
end 13'h3ec:    begin Red = 8'h71;    Green = 8'h78;    Blue = 8'h5b;
end 13'h3ed:    begin Red = 8'h7c;    Green = 8'h8c;    Blue = 8'h40;
end 13'h3ee:    begin Red = 8'hd2;    Green = 8'hc7;    Blue = 8'hca;
end 13'h3ef:    begin Red = 8'hb8;    Green = 8'hc2;    Blue = 8'hbe;
end 13'h3f0:    begin Red = 8'hb5;    Green = 8'hc1;    Blue = 8'hbb;
end 13'h3f1:    begin Red = 8'hcf;    Green = 8'hce;    Blue = 8'hd3;
end 13'h3f2:    begin Red = 8'h7d;    Green = 8'h90;    Blue = 8'h51;
end 13'h3f3:    begin Red = 8'h8b;    Green = 8'h90;    Blue = 8'h78;
end 13'h3f4:    begin Red = 8'h7f;    Green = 8'h85;    Blue = 8'h79;
end 13'h3f5:    begin Red = 8'ha8;    Green = 8'haf;    Blue = 8'hac;
end 13'h3f6:    begin Red = 8'hac;    Green = 8'hb3;    Blue = 8'haf;
end 13'h3f7:    begin Red = 8'hab;    Green = 8'hb0;    Blue = 8'hab;
end 13'h3f8:    begin Red = 8'h6e;    Green = 8'h6c;    Blue = 8'h62;
end 13'h3f9:    begin Red = 8'h70;    Green = 8'h69;    Blue = 8'h5f;
end 13'h3fa:    begin Red = 8'h88;    Green = 8'h91;    Blue = 8'h5a;
end 13'h3fb:    begin Red = 8'h82;    Green = 8'h81;    Blue = 8'h5b;
end 13'h3fc:    begin Red = 8'hb0;    Green = 8'hab;    Blue = 8'h55;
end 13'h3fd:    begin Red = 8'ha1;    Green = 8'h9f;    Blue = 8'h4a;
end 13'h3fe:    begin Red = 8'ha3;    Green = 8'h9a;    Blue = 8'h52;
end 13'h3ff:    begin Red = 8'h98;    Green = 8'h9e;    Blue = 8'h51;
end 13'h400:    begin Red = 8'hbe;    Green = 8'hc1;    Blue = 8'h4d;
end 13'h401:    begin Red = 8'h9e;    Green = 8'ha7;    Blue = 8'h50;
end 13'h402:    begin Red = 8'hb5;    Green = 8'ha9;    Blue = 8'h44;
end 13'h403:    begin Red = 8'hd2;    Green = 8'hbd;    Blue = 8'h99;
end 13'h404:    begin Red = 8'hba;    Green = 8'ha1;    Blue = 8'h8a;
end 13'h405:    begin Red = 8'hbd;    Green = 8'ha6;    Blue = 8'h8c;
end 13'h406:    begin Red = 8'h6b;    Green = 8'h73;    Blue = 8'h49;
end 13'h407:    begin Red = 8'h74;    Green = 8'h80;    Blue = 8'h4f;
end 13'h408:    begin Red = 8'h82;    Green = 8'h98;    Blue = 8'h40;
end 13'h409:    begin Red = 8'h9e;    Green = 8'hb2;    Blue = 8'h98;
end 13'h40a:    begin Red = 8'h8d;    Green = 8'haf;    Blue = 8'h8f;
end 13'h40b:    begin Red = 8'hd3;    Green = 8'hd2;    Blue = 8'hce;
end 13'h40c:    begin Red = 8'hd4;    Green = 8'hd5;    Blue = 8'hca;
end 13'h40d:    begin Red = 8'h7c;    Green = 8'h94;    Blue = 8'h7d;
end 13'h40e:    begin Red = 8'hdc;    Green = 8'hdd;    Blue = 8'he1;
end 13'h40f:    begin Red = 8'hd2;    Green = 8'hd2;    Blue = 8'hca;
end 13'h410:    begin Red = 8'h97;    Green = 8'haf;    Blue = 8'h94;
end 13'h411:    begin Red = 8'hc3;    Green = 8'hc3;    Blue = 8'hbf;
end 13'h412:    begin Red = 8'he0;    Green = 8'hdc;    Blue = 8'hdf;
end 13'h413:    begin Red = 8'h6d;    Green = 8'h7c;    Blue = 8'h67;
end 13'h414:    begin Red = 8'hcc;    Green = 8'hc8;    Blue = 8'haa;
end 13'h415:    begin Red = 8'hc2;    Green = 8'hc0;    Blue = 8'ha2;
end 13'h416:    begin Red = 8'h96;    Green = 8'h98;    Blue = 8'h83;
end 13'h417:    begin Red = 8'h73;    Green = 8'h79;    Blue = 8'h4c;
end 13'h418:    begin Red = 8'h8c;    Green = 8'h9b;    Blue = 8'h5a;
end 13'h419:    begin Red = 8'h8d;    Green = 8'h9d;    Blue = 8'h56;
end 13'h41a:    begin Red = 8'hbb;    Green = 8'h91;    Blue = 8'h70;
end 13'h41b:    begin Red = 8'hb3;    Green = 8'h8c;    Blue = 8'h6a;
end 13'h41c:    begin Red = 8'h9b;    Green = 8'ha3;    Blue = 8'h5c;
end 13'h41d:    begin Red = 8'h8c;    Green = 8'h88;    Blue = 8'h78;
end 13'h41e:    begin Red = 8'h8a;    Green = 8'h88;    Blue = 8'h7c;
end 13'h41f:    begin Red = 8'h8a;    Green = 8'h92;    Blue = 8'h89;
end 13'h420:    begin Red = 8'h94;    Green = 8'h78;    Blue = 8'h5e;
end 13'h421:    begin Red = 8'ha3;    Green = 8'h87;    Blue = 8'h6c;
end 13'h422:    begin Red = 8'ha5;    Green = 8'h82;    Blue = 8'h65;
end 13'h423:    begin Red = 8'h6d;    Green = 8'h66;    Blue = 8'h67;
end 13'h424:    begin Red = 8'h67;    Green = 8'h69;    Blue = 8'h5c;
end 13'h425:    begin Red = 8'h65;    Green = 8'h64;    Blue = 8'h5a;
end 13'h426:    begin Red = 8'h9f;    Green = 8'hb3;    Blue = 8'h4b;
end 13'h427:    begin Red = 8'h7b;    Green = 8'h86;    Blue = 8'h57;
end 13'h428:    begin Red = 8'h7e;    Green = 8'h78;    Blue = 8'h61;
end 13'h429:    begin Red = 8'h8c;    Green = 8'h7a;    Blue = 8'h5a;
end 13'h42a:    begin Red = 8'h8c;    Green = 8'h82;    Blue = 8'h58;
end 13'h42b:    begin Red = 8'hb6;    Green = 8'haf;    Blue = 8'h50;
end 13'h42c:    begin Red = 8'hae;    Green = 8'haa;    Blue = 8'h4c;
end 13'h42d:    begin Red = 8'haa;    Green = 8'ha1;    Blue = 8'h4e;
end 13'h42e:    begin Red = 8'h9f;    Green = 8'h9b;    Blue = 8'h5a;
end 13'h42f:    begin Red = 8'hce;    Green = 8'hc5;    Blue = 8'h59;
end 13'h430:    begin Red = 8'h9b;    Green = 8'h9b;    Blue = 8'h51;
end 13'h431:    begin Red = 8'ha7;    Green = 8'h9f;    Blue = 8'h51;
end 13'h432:    begin Red = 8'h50;    Green = 8'h6f;    Blue = 8'h88;
end 13'h433:    begin Red = 8'h51;    Green = 8'h74;    Blue = 8'h7b;
end 13'h434:    begin Red = 8'h51;    Green = 8'h73;    Blue = 8'h80;
end 13'h435:    begin Red = 8'h64;    Green = 8'h78;    Blue = 8'h79;
end 13'h436:    begin Red = 8'he1;    Green = 8'hc5;    Blue = 8'ha7;
end 13'h437:    begin Red = 8'hd6;    Green = 8'hbb;    Blue = 8'ha3;
end 13'h438:    begin Red = 8'h80;    Green = 8'h6b;    Blue = 8'h55;
end 13'h439:    begin Red = 8'hc5;    Green = 8'had;    Blue = 8'h97;
end 13'h43a:    begin Red = 8'hfd;    Green = 8'hff;    Blue = 8'hea;
end 13'h43b:    begin Red = 8'hfb;    Green = 8'hf6;    Blue = 8'hd9;
end 13'h43c:    begin Red = 8'ha2;    Green = 8'hb9;    Blue = 8'h5a;
end 13'h43d:    begin Red = 8'h94;    Green = 8'ha7;    Blue = 8'h46;
end 13'h43e:    begin Red = 8'hff;    Green = 8'hea;    Blue = 8'hd9;
end 13'h43f:    begin Red = 8'h96;    Green = 8'hb6;    Blue = 8'ha3;
end 13'h440:    begin Red = 8'h99;    Green = 8'hbb;    Blue = 8'h9e;
end 13'h441:    begin Red = 8'hed;    Green = 8'hf5;    Blue = 8'hf1;
end 13'h442:    begin Red = 8'he2;    Green = 8'hec;    Blue = 8'hf2;
end 13'h443:    begin Red = 8'he7;    Green = 8'he3;    Blue = 8'he0;
end 13'h444:    begin Red = 8'hdd;    Green = 8'he2;    Blue = 8'hd6;
end 13'h445:    begin Red = 8'hde;    Green = 8'he4;    Blue = 8'he5;
end 13'h446:    begin Red = 8'he1;    Green = 8'he2;    Blue = 8'hdd;
end 13'h447:    begin Red = 8'he2;    Green = 8'hda;    Blue = 8'he3;
end 13'h448:    begin Red = 8'hf0;    Green = 8'hf0;    Blue = 8'hf0;
end 13'h449:    begin Red = 8'hd8;    Green = 8'he0;    Blue = 8'hd7;
end 13'h44a:    begin Red = 8'hd4;    Green = 8'hd1;    Blue = 8'hc7;
end 13'h44b:    begin Red = 8'hde;    Green = 8'hdf;    Blue = 8'he9;
end 13'h44c:    begin Red = 8'h93;    Green = 8'hb1;    Blue = 8'h92;
end 13'h44d:    begin Red = 8'he8;    Green = 8'he7;    Blue = 8'hec;
end 13'h44e:    begin Red = 8'hd9;    Green = 8'he2;    Blue = 8'hda;
end 13'h44f:    begin Red = 8'hd1;    Green = 8'hd4;    Blue = 8'hc8;
end 13'h450:    begin Red = 8'hea;    Green = 8'hde;    Blue = 8'he0;
end 13'h451:    begin Red = 8'he2;    Green = 8'hdb;    Blue = 8'hea;
end 13'h452:    begin Red = 8'hd9;    Green = 8'hd2;    Blue = 8'hca;
end 13'h453:    begin Red = 8'h65;    Green = 8'h78;    Blue = 8'h65;
end 13'h454:    begin Red = 8'h65;    Green = 8'h82;    Blue = 8'h64;
end 13'h455:    begin Red = 8'hc1;    Green = 8'hc7;    Blue = 8'hc0;
end 13'h456:    begin Red = 8'hc3;    Green = 8'hc7;    Blue = 8'hb9;
end 13'h457:    begin Red = 8'h5d;    Green = 8'h6e;    Blue = 8'h5c;
end 13'h458:    begin Red = 8'h72;    Green = 8'h86;    Blue = 8'h6f;
end 13'h459:    begin Red = 8'h6e;    Green = 8'h88;    Blue = 8'h70;
end 13'h45a:    begin Red = 8'hca;    Green = 8'hd2;    Blue = 8'hcb;
end 13'h45b:    begin Red = 8'h59;    Green = 8'h70;    Blue = 8'h5e;
end 13'h45c:    begin Red = 8'h59;    Green = 8'h6d;    Blue = 8'h5a;
end 13'h45d:    begin Red = 8'hd6;    Green = 8'hd2;    Blue = 8'hd5;
end 13'h45e:    begin Red = 8'h5a;    Green = 8'h72;    Blue = 8'h7b;
end 13'h45f:    begin Red = 8'hbf;    Green = 8'hc0;    Blue = 8'ha5;
end 13'h460:    begin Red = 8'h98;    Green = 8'h9d;    Blue = 8'h95;
end 13'h461:    begin Red = 8'h9e;    Green = 8'h9c;    Blue = 8'h93;
end 13'h462:    begin Red = 8'h76;    Green = 8'h7f;    Blue = 8'h51;
end 13'h463:    begin Red = 8'hca;    Green = 8'h98;    Blue = 8'h7f;
end 13'h464:    begin Red = 8'hc4;    Green = 8'h96;    Blue = 8'h6e;
end 13'h465:    begin Red = 8'h7e;    Green = 8'h7d;    Blue = 8'h4c;
end 13'h466:    begin Red = 8'h80;    Green = 8'h7f;    Blue = 8'h51;
end 13'h467:    begin Red = 8'h99;    Green = 8'h95;    Blue = 8'h93;
end 13'h468:    begin Red = 8'h88;    Green = 8'h82;    Blue = 8'h88;
end 13'h469:    begin Red = 8'h88;    Green = 8'h83;    Blue = 8'h84;
end 13'h46a:    begin Red = 8'h84;    Green = 8'h88;    Blue = 8'h8b;
end 13'h46b:    begin Red = 8'ha3;    Green = 8'h8a;    Blue = 8'h63;
end 13'h46c:    begin Red = 8'ha0;    Green = 8'h82;    Blue = 8'h63;
end 13'h46d:    begin Red = 8'hac;    Green = 8'hc3;    Blue = 8'h4c;
end 13'h46e:    begin Red = 8'hb5;    Green = 8'hcf;    Blue = 8'h44;
end 13'h46f:    begin Red = 8'h87;    Green = 8'h95;    Blue = 8'h52;
end 13'h470:    begin Red = 8'h9c;    Green = 8'hb1;    Blue = 8'h45;
end 13'h471:    begin Red = 8'h80;    Green = 8'h89;    Blue = 8'h61;
end 13'h472:    begin Red = 8'h9e;    Green = 8'hb4;    Blue = 8'h41;
end 13'h473:    begin Red = 8'h83;    Green = 8'h8c;    Blue = 8'h5a;
end 13'h474:    begin Red = 8'h94;    Green = 8'h93;    Blue = 8'h51;
end 13'h475:    begin Red = 8'h8e;    Green = 8'h7f;    Blue = 8'h5d;
end 13'h476:    begin Red = 8'h9d;    Green = 8'ha3;    Blue = 8'h57;
end 13'h477:    begin Red = 8'hc7;    Green = 8'hbf;    Blue = 8'h57;
end 13'h478:    begin Red = 8'hc4;    Green = 8'hbd;    Blue = 8'h60;
end 13'h479:    begin Red = 8'hb3;    Green = 8'h9d;    Blue = 8'h92;
end 13'h47a:    begin Red = 8'haa;    Green = 8'ha3;    Blue = 8'h8c;
end 13'h47b:    begin Red = 8'h4a;    Green = 8'h70;    Blue = 8'h7d;
end 13'h47c:    begin Red = 8'h95;    Green = 8'h86;    Blue = 8'h6c;
end 13'h47d:    begin Red = 8'h94;    Green = 8'h84;    Blue = 8'h71;
end 13'h47e:    begin Red = 8'h8b;    Green = 8'h7e;    Blue = 8'h61;
end 13'h47f:    begin Red = 8'h87;    Green = 8'h8c;    Blue = 8'h55;
end 13'h480:    begin Red = 8'h8d;    Green = 8'h93;    Blue = 8'h5b;
end 13'h481:    begin Red = 8'h5c;    Green = 8'h61;    Blue = 8'h47;
end 13'h482:    begin Red = 8'h55;    Green = 8'h5d;    Blue = 8'h3b;
end 13'h483:    begin Red = 8'h5b;    Green = 8'h64;    Blue = 8'h36;
end 13'h484:    begin Red = 8'h67;    Green = 8'h73;    Blue = 8'h47;
end 13'h485:    begin Red = 8'h6c;    Green = 8'h66;    Blue = 8'h5a;
end 13'h486:    begin Red = 8'ha0;    Green = 8'hb1;    Blue = 8'had;
end 13'h487:    begin Red = 8'h90;    Green = 8'hbd;    Blue = 8'ha0;
end 13'h488:    begin Red = 8'hb1;    Green = 8'ha3;    Blue = 8'h8c;
end 13'h489:    begin Red = 8'he8;    Green = 8'hdd;    Blue = 8'hdc;
end 13'h48a:    begin Red = 8'h96;    Green = 8'hb7;    Blue = 8'h94;
end 13'h48b:    begin Red = 8'ha6;    Green = 8'ha7;    Blue = 8'ha3;
end 13'h48c:    begin Red = 8'ha8;    Green = 8'ha8;    Blue = 8'ha7;
end 13'h48d:    begin Red = 8'haf;    Green = 8'hae;    Blue = 8'hab;
end 13'h48e:    begin Red = 8'hcb;    Green = 8'hd2;    Blue = 8'hc5;
end 13'h48f:    begin Red = 8'hac;    Green = 8'ha7;    Blue = 8'hab;
end 13'h490:    begin Red = 8'ha3;    Green = 8'ha8;    Blue = 8'ha2;
end 13'h491:    begin Red = 8'hba;    Green = 8'ha9;    Blue = 8'ha7;
end 13'h492:    begin Red = 8'he8;    Green = 8'he2;    Blue = 8'he9;
end 13'h493:    begin Red = 8'hcf;    Green = 8'hd1;    Blue = 8'hcd;
end 13'h494:    begin Red = 8'he1;    Green = 8'hd8;    Blue = 8'hd3;
end 13'h495:    begin Red = 8'hbc;    Green = 8'hbe;    Blue = 8'hb9;
end 13'h496:    begin Red = 8'hc2;    Green = 8'hbe;    Blue = 8'hb9;
end 13'h497:    begin Red = 8'hcb;    Green = 8'hce;    Blue = 8'hcf;
end 13'h498:    begin Red = 8'hcd;    Green = 8'hcb;    Blue = 8'hcc;
end 13'h499:    begin Red = 8'hbf;    Green = 8'hc1;    Blue = 8'hb7;
end 13'h49a:    begin Red = 8'hc3;    Green = 8'hbf;    Blue = 8'hbd;
end 13'h49b:    begin Red = 8'hcc;    Green = 8'hce;    Blue = 8'hcb;
end 13'h49c:    begin Red = 8'hca;    Green = 8'hcb;    Blue = 8'hce;
end 13'h49d:    begin Red = 8'hc9;    Green = 8'hce;    Blue = 8'hc6;
end 13'h49e:    begin Red = 8'hc7;    Green = 8'hbf;    Blue = 8'hc0;
end 13'h49f:    begin Red = 8'h56;    Green = 8'h72;    Blue = 8'h61;
end 13'h4a0:    begin Red = 8'h6c;    Green = 8'h7d;    Blue = 8'h6f;
end 13'h4a1:    begin Red = 8'h8d;    Green = 8'h97;    Blue = 8'h78;
end 13'h4a2:    begin Red = 8'hc3;    Green = 8'hc2;    Blue = 8'hac;
end 13'h4a3:    begin Red = 8'h71;    Green = 8'h7f;    Blue = 8'h46;
end 13'h4a4:    begin Red = 8'h60;    Green = 8'h65;    Blue = 8'h44;
end 13'h4a5:    begin Red = 8'h79;    Green = 8'h8a;    Blue = 8'h53;
end 13'h4a6:    begin Red = 8'h68;    Green = 8'h58;    Blue = 8'h5f;
end 13'h4a7:    begin Red = 8'h81;    Green = 8'h8c;    Blue = 8'h5f;
end 13'h4a8:    begin Red = 8'h9e;    Green = 8'hb3;    Blue = 8'h47;
end 13'h4a9:    begin Red = 8'h96;    Green = 8'hb4;    Blue = 8'h3f;
end 13'h4aa:    begin Red = 8'h90;    Green = 8'h76;    Blue = 8'h57;
end 13'h4ab:    begin Red = 8'hac;    Green = 8'h8b;    Blue = 8'h66;
end 13'h4ac:    begin Red = 8'h9b;    Green = 8'had;    Blue = 8'h52;
end 13'h4ad:    begin Red = 8'h7b;    Green = 8'h8d;    Blue = 8'h57;
end 13'h4ae:    begin Red = 8'h98;    Green = 8'had;    Blue = 8'h46;
end 13'h4af:    begin Red = 8'ha0;    Green = 8'hb6;    Blue = 8'h44;
end 13'h4b0:    begin Red = 8'h98;    Green = 8'hac;    Blue = 8'h4c;
end 13'h4b1:    begin Red = 8'had;    Green = 8'hb7;    Blue = 8'h37;
end 13'h4b2:    begin Red = 8'h55;    Green = 8'h77;    Blue = 8'h7c;
end 13'h4b3:    begin Red = 8'hae;    Green = 8'h9d;    Blue = 8'h5e;
end 13'h4b4:    begin Red = 8'h9e;    Green = 8'ha4;    Blue = 8'h54;
end 13'h4b5:    begin Red = 8'ha3;    Green = 8'h9e;    Blue = 8'h56;
end 13'h4b6:    begin Red = 8'hb3;    Green = 8'ha2;    Blue = 8'h93;
end 13'h4b7:    begin Red = 8'h4e;    Green = 8'h74;    Blue = 8'h77;
end 13'h4b8:    begin Red = 8'h95;    Green = 8'h88;    Blue = 8'h74;
end 13'h4b9:    begin Red = 8'hd7;    Green = 8'hbf;    Blue = 8'ha1;
end 13'h4ba:    begin Red = 8'ha6;    Green = 8'h91;    Blue = 8'h7d;
end 13'h4bb:    begin Red = 8'h79;    Green = 8'h82;    Blue = 8'h52;
end 13'h4bc:    begin Red = 8'h60;    Green = 8'h61;    Blue = 8'h46;
end 13'h4bd:    begin Red = 8'h77;    Green = 8'h84;    Blue = 8'h4a;
end 13'h4be:    begin Red = 8'h6a;    Green = 8'h6d;    Blue = 8'h62;
end 13'h4bf:    begin Red = 8'h6e;    Green = 8'h72;    Blue = 8'h5a;
end 13'h4c0:    begin Red = 8'hb0;    Green = 8'hc9;    Blue = 8'h47;
end 13'h4c1:    begin Red = 8'haf;    Green = 8'hc8;    Blue = 8'h34;
end 13'h4c2:    begin Red = 8'hb4;    Green = 8'ha0;    Blue = 8'h85;
end 13'h4c3:    begin Red = 8'haf;    Green = 8'ha3;    Blue = 8'h89;
end 13'h4c4:    begin Red = 8'haf;    Green = 8'ha0;    Blue = 8'h87;
end 13'h4c5:    begin Red = 8'h9a;    Green = 8'ha3;    Blue = 8'h9c;
end 13'h4c6:    begin Red = 8'hab;    Green = 8'ha2;    Blue = 8'ha8;
end 13'h4c7:    begin Red = 8'h9e;    Green = 8'ha3;    Blue = 8'h9d;
end 13'h4c8:    begin Red = 8'h9b;    Green = 8'hbc;    Blue = 8'h9b;
end 13'h4c9:    begin Red = 8'h9c;    Green = 8'ha1;    Blue = 8'h9e;
end 13'h4ca:    begin Red = 8'ha2;    Green = 8'h9e;    Blue = 8'h9b;
end 13'h4cb:    begin Red = 8'hac;    Green = 8'ha5;    Blue = 8'ha7;
end 13'h4cc:    begin Red = 8'h7c;    Green = 8'h99;    Blue = 8'h7f;
end 13'h4cd:    begin Red = 8'ha4;    Green = 8'ha2;    Blue = 8'ha9;
end 13'h4ce:    begin Red = 8'ha1;    Green = 8'h9b;    Blue = 8'ha2;
end 13'h4cf:    begin Red = 8'ha1;    Green = 8'h9c;    Blue = 8'ha7;
end 13'h4d0:    begin Red = 8'h9f;    Green = 8'ha2;    Blue = 8'ha3;
end 13'h4d1:    begin Red = 8'h84;    Green = 8'h92;    Blue = 8'h85;
end 13'h4d2:    begin Red = 8'h8e;    Green = 8'h98;    Blue = 8'h93;
end 13'h4d3:    begin Red = 8'ha1;    Green = 8'ha0;    Blue = 8'ha2;
end 13'h4d4:    begin Red = 8'h95;    Green = 8'h97;    Blue = 8'h93;
end 13'h4d5:    begin Red = 8'he9;    Green = 8'he2;    Blue = 8'hee;
end 13'h4d6:    begin Red = 8'hd2;    Green = 8'hcb;    Blue = 8'hc9;
end 13'h4d7:    begin Red = 8'h88;    Green = 8'h90;    Blue = 8'h7a;
end 13'h4d8:    begin Red = 8'hcf;    Green = 8'hca;    Blue = 8'hcf;
end 13'h4d9:    begin Red = 8'h75;    Green = 8'h7f;    Blue = 8'h78;
end 13'h4da:    begin Red = 8'h69;    Green = 8'h80;    Blue = 8'h6e;
end 13'h4db:    begin Red = 8'h8a;    Green = 8'h99;    Blue = 8'h88;
end 13'h4dc:    begin Red = 8'hca;    Green = 8'hc4;    Blue = 8'ha7;
end 13'h4dd:    begin Red = 8'hb9;    Green = 8'hbb;    Blue = 8'ha3;
end 13'h4de:    begin Red = 8'h94;    Green = 8'h98;    Blue = 8'h86;
end 13'h4df:    begin Red = 8'h62;    Green = 8'h72;    Blue = 8'h43;
end 13'h4e0:    begin Red = 8'h6d;    Green = 8'h7d;    Blue = 8'h46;
end 13'h4e1:    begin Red = 8'h5a;    Green = 8'h5f;    Blue = 8'h4a;
end 13'h4e2:    begin Red = 8'h54;    Green = 8'h60;    Blue = 8'h41;
end 13'h4e3:    begin Red = 8'h65;    Green = 8'h63;    Blue = 8'h44;
end 13'h4e4:    begin Red = 8'h72;    Green = 8'h6e;    Blue = 8'h5e;
end 13'h4e5:    begin Red = 8'h7c;    Green = 8'h8c;    Blue = 8'h5f;
end 13'h4e6:    begin Red = 8'hab;    Green = 8'hc3;    Blue = 8'h48;
end 13'h4e7:    begin Red = 8'ha2;    Green = 8'hba;    Blue = 8'h3c;
end 13'h4e8:    begin Red = 8'h83;    Green = 8'h90;    Blue = 8'h52;
end 13'h4e9:    begin Red = 8'h7f;    Green = 8'h8a;    Blue = 8'h5b;
end 13'h4ea:    begin Red = 8'h82;    Green = 8'h8c;    Blue = 8'h64;
end 13'h4eb:    begin Red = 8'h7f;    Green = 8'h8b;    Blue = 8'h55;
end 13'h4ec:    begin Red = 8'ha9;    Green = 8'hc1;    Blue = 8'h42;
end 13'h4ed:    begin Red = 8'ha1;    Green = 8'hb8;    Blue = 8'h3f;
end 13'h4ee:    begin Red = 8'h78;    Green = 8'h83;    Blue = 8'h59;
end 13'h4ef:    begin Red = 8'hb3;    Green = 8'hc1;    Blue = 8'h4b;
end 13'h4f0:    begin Red = 8'hb2;    Green = 8'hce;    Blue = 8'h38;
end 13'h4f1:    begin Red = 8'h64;    Green = 8'h81;    Blue = 8'h97;
end 13'h4f2:    begin Red = 8'h50;    Green = 8'h6f;    Blue = 8'h7b;
end 13'h4f3:    begin Red = 8'h46;    Green = 8'h6c;    Blue = 8'h7e;
end 13'h4f4:    begin Red = 8'h52;    Green = 8'h6c;    Blue = 8'h78;
end 13'h4f5:    begin Red = 8'h3e;    Green = 8'h6b;    Blue = 8'h82;
end 13'h4f6:    begin Red = 8'hb5;    Green = 8'h9d;    Blue = 8'h8a;
end 13'h4f7:    begin Red = 8'ha0;    Green = 8'ha3;    Blue = 8'h46;
end 13'h4f8:    begin Red = 8'h9e;    Green = 8'ha1;    Blue = 8'h49;
end 13'h4f9:    begin Red = 8'hac;    Green = 8'ha2;    Blue = 8'h94;
end 13'h4fa:    begin Red = 8'h48;    Green = 8'h6a;    Blue = 8'h79;
end 13'h4fb:    begin Red = 8'h43;    Green = 8'h65;    Blue = 8'h75;
end 13'h4fc:    begin Red = 8'h47;    Green = 8'h72;    Blue = 8'h7a;
end 13'h4fd:    begin Red = 8'h53;    Green = 8'h6b;    Blue = 8'h81;
end 13'h4fe:    begin Red = 8'h7e;    Green = 8'h68;    Blue = 8'h5d;
end 13'h4ff:    begin Red = 8'h7d;    Green = 8'h69;    Blue = 8'h59;
end 13'h500:    begin Red = 8'h60;    Green = 8'h7e;    Blue = 8'h42;
end 13'h501:    begin Red = 8'h75;    Green = 8'h90;    Blue = 8'h47;
end 13'h502:    begin Red = 8'h6c;    Green = 8'h7b;    Blue = 8'h48;
end 13'h503:    begin Red = 8'h5b;    Green = 8'h61;    Blue = 8'h41;
end 13'h504:    begin Red = 8'h78;    Green = 8'h84;    Blue = 8'h55;
end 13'h505:    begin Red = 8'h75;    Green = 8'h81;    Blue = 8'h4a;
end 13'h506:    begin Red = 8'h74;    Green = 8'h81;    Blue = 8'h43;
end 13'h507:    begin Red = 8'h6b;    Green = 8'h6d;    Blue = 8'h5d;
end 13'h508:    begin Red = 8'h62;    Green = 8'h5a;    Blue = 8'h5b;
end 13'h509:    begin Red = 8'h76;    Green = 8'h89;    Blue = 8'h5a;
end 13'h50a:    begin Red = 8'ha1;    Green = 8'hb4;    Blue = 8'h3d;
end 13'h50b:    begin Red = 8'h91;    Green = 8'haf;    Blue = 8'h3c;
end 13'h50c:    begin Red = 8'ha5;    Green = 8'hc7;    Blue = 8'h3c;
end 13'h50d:    begin Red = 8'h9a;    Green = 8'hc2;    Blue = 8'h36;
end 13'h50e:    begin Red = 8'h8e;    Green = 8'hb0;    Blue = 8'h98;
end 13'h50f:    begin Red = 8'h86;    Green = 8'hbb;    Blue = 8'h94;
end 13'h510:    begin Red = 8'h9b;    Green = 8'h98;    Blue = 8'haa;
end 13'h511:    begin Red = 8'h99;    Green = 8'h9a;    Blue = 8'ha8;
end 13'h512:    begin Red = 8'h6e;    Green = 8'h8b;    Blue = 8'h76;
end 13'h513:    begin Red = 8'h95;    Green = 8'hb7;    Blue = 8'ha0;
end 13'h514:    begin Red = 8'h90;    Green = 8'hb3;    Blue = 8'h98;
end 13'h515:    begin Red = 8'h8b;    Green = 8'hb3;    Blue = 8'h94;
end 13'h516:    begin Red = 8'h8c;    Green = 8'h9e;    Blue = 8'h9c;
end 13'h517:    begin Red = 8'h6d;    Green = 8'h84;    Blue = 8'h76;
end 13'h518:    begin Red = 8'h8a;    Green = 8'hac;    Blue = 8'h96;
end 13'h519:    begin Red = 8'h90;    Green = 8'hb0;    Blue = 8'h9b;
end 13'h51a:    begin Red = 8'h91;    Green = 8'hae;    Blue = 8'h99;
end 13'h51b:    begin Red = 8'ha4;    Green = 8'hb4;    Blue = 8'h9e;
end 13'h51c:    begin Red = 8'h99;    Green = 8'hbe;    Blue = 8'h99;
end 13'h51d:    begin Red = 8'ha0;    Green = 8'h98;    Blue = 8'h9f;
end 13'h51e:    begin Red = 8'h9f;    Green = 8'hb5;    Blue = 8'ha3;
end 13'h51f:    begin Red = 8'haa;    Green = 8'h9e;    Blue = 8'ha3;
end 13'h520:    begin Red = 8'h7a;    Green = 8'h90;    Blue = 8'h72;
end 13'h521:    begin Red = 8'ha8;    Green = 8'ha0;    Blue = 8'ha9;
end 13'h522:    begin Red = 8'ha2;    Green = 8'ha2;    Blue = 8'ha0;
end 13'h523:    begin Red = 8'ha3;    Green = 8'h9d;    Blue = 8'ha3;
end 13'h524:    begin Red = 8'h9b;    Green = 8'h9b;    Blue = 8'h9d;
end 13'h525:    begin Red = 8'h75;    Green = 8'h8e;    Blue = 8'h75;
end 13'h526:    begin Red = 8'hed;    Green = 8'he0;    Blue = 8'he9;
end 13'h527:    begin Red = 8'h9b;    Green = 8'h98;    Blue = 8'h98;
end 13'h528:    begin Red = 8'h9e;    Green = 8'h98;    Blue = 8'ha3;
end 13'h529:    begin Red = 8'he3;    Green = 8'hd6;    Blue = 8'hda;
end 13'h52a:    begin Red = 8'hdb;    Green = 8'hd9;    Blue = 8'hd2;
end 13'h52b:    begin Red = 8'hde;    Green = 8'hd6;    Blue = 8'hde;
end 13'h52c:    begin Red = 8'hd6;    Green = 8'hca;    Blue = 8'hca;
end 13'h52d:    begin Red = 8'h6e;    Green = 8'h78;    Blue = 8'h71;
end 13'h52e:    begin Red = 8'hdf;    Green = 8'hde;    Blue = 8'hed;
end 13'h52f:    begin Red = 8'hcf;    Green = 8'hca;    Blue = 8'hca;
end 13'h530:    begin Red = 8'h75;    Green = 8'h98;    Blue = 8'h82;
end 13'h531:    begin Red = 8'h71;    Green = 8'h8e;    Blue = 8'h80;
end 13'h532:    begin Red = 8'h42;    Green = 8'h67;    Blue = 8'h7c;
end 13'h533:    begin Red = 8'h47;    Green = 8'h6e;    Blue = 8'h79;
end 13'h534:    begin Red = 8'h4d;    Green = 8'h6e;    Blue = 8'h80;
end 13'h535:    begin Red = 8'hbe;    Green = 8'hc7;    Blue = 8'had;
end 13'h536:    begin Red = 8'h5d;    Green = 8'h6b;    Blue = 8'h3a;
end 13'h537:    begin Red = 8'h8d;    Green = 8'h9c;    Blue = 8'h46;
end 13'h538:    begin Red = 8'h72;    Green = 8'h7c;    Blue = 8'h47;
end 13'h539:    begin Red = 8'h74;    Green = 8'h89;    Blue = 8'h4c;
end 13'h53a:    begin Red = 8'h73;    Green = 8'h84;    Blue = 8'h48;
end 13'h53b:    begin Red = 8'h71;    Green = 8'h6e;    Blue = 8'h65;
end 13'h53c:    begin Red = 8'h6c;    Green = 8'h69;    Blue = 8'h60;
end 13'h53d:    begin Red = 8'h6e;    Green = 8'h88;    Blue = 8'h4a;
end 13'h53e:    begin Red = 8'h6c;    Green = 8'h82;    Blue = 8'h51;
end 13'h53f:    begin Red = 8'h8c;    Green = 8'hac;    Blue = 8'h3c;
end 13'h540:    begin Red = 8'h9e;    Green = 8'hc5;    Blue = 8'h3e;
end 13'h541:    begin Red = 8'h9e;    Green = 8'hc7;    Blue = 8'h37;
end 13'h542:    begin Red = 8'hae;    Green = 8'hc6;    Blue = 8'h48;
end 13'h543:    begin Red = 8'h9a;    Green = 8'haf;    Blue = 8'h42;
end 13'h544:    begin Red = 8'h53;    Green = 8'h51;    Blue = 8'h4b;
end 13'h545:    begin Red = 8'hfa;    Green = 8'he2;    Blue = 8'hb7;
end 13'h546:    begin Red = 8'hd9;    Green = 8'hca;    Blue = 8'ha4;
end 13'h547:    begin Red = 8'hec;    Green = 8'hcd;    Blue = 8'hb4;
end 13'h548:    begin Red = 8'hb8;    Green = 8'h9d;    Blue = 8'h88;
end 13'h549:    begin Red = 8'hc9;    Green = 8'hbd;    Blue = 8'h9b;
end 13'h54a:    begin Red = 8'hda;    Green = 8'hc8;    Blue = 8'ha7;
end 13'h54b:    begin Red = 8'hdf;    Green = 8'hc9;    Blue = 8'haa;
end 13'h54c:    begin Red = 8'hfb;    Green = 8'he5;    Blue = 8'hce;
end 13'h54d:    begin Red = 8'hdf;    Green = 8'hc3;    Blue = 8'ha5;
end 13'h54e:    begin Red = 8'h90;    Green = 8'h7a;    Blue = 8'h69;
end 13'h54f:    begin Red = 8'hc6;    Green = 8'haf;    Blue = 8'h9e;
end 13'h550:    begin Red = 8'ha9;    Green = 8'h90;    Blue = 8'h78;
end 13'h551:    begin Red = 8'h5f;    Green = 8'h65;    Blue = 8'h48;
end 13'h552:    begin Red = 8'h5a;    Green = 8'h60;    Blue = 8'h3d;
end 13'h553:    begin Red = 8'hc4;    Green = 8'hac;    Blue = 8'h8e;
end 13'h554:    begin Red = 8'hc4;    Green = 8'haf;    Blue = 8'h8c;
end 13'h555:    begin Red = 8'he5;    Green = 8'hce;    Blue = 8'haf;
end 13'h556:    begin Red = 8'he0;    Green = 8'hc9;    Blue = 8'hb1;
end 13'h557:    begin Red = 8'he3;    Green = 8'hc9;    Blue = 8'ha5;
end 13'h558:    begin Red = 8'he2;    Green = 8'hca;    Blue = 8'ha2;
end 13'h559:    begin Red = 8'hec;    Green = 8'hd5;    Blue = 8'hb2;
end 13'h55a:    begin Red = 8'hc8;    Green = 8'hb8;    Blue = 8'h9b;
end 13'h55b:    begin Red = 8'hdf;    Green = 8'hca;    Blue = 8'ha4;
end 13'h55c:    begin Red = 8'he2;    Green = 8'hcc;    Blue = 8'ha7;
end 13'h55d:    begin Red = 8'h96;    Green = 8'hb7;    Blue = 8'h9b;
end 13'h55e:    begin Red = 8'h9e;    Green = 8'hb1;    Blue = 8'ha4;
end 13'h55f:    begin Red = 8'h9b;    Green = 8'h9e;    Blue = 8'h98;
end 13'h560:    begin Red = 8'ha0;    Green = 8'h97;    Blue = 8'h9a;
end 13'h561:    begin Red = 8'h9e;    Green = 8'h9e;    Blue = 8'h9c;
end 13'h562:    begin Red = 8'h7f;    Green = 8'h93;    Blue = 8'h81;
end 13'h563:    begin Red = 8'h9a;    Green = 8'h9b;    Blue = 8'h96;
end 13'h564:    begin Red = 8'ha7;    Green = 8'h9f;    Blue = 8'ha0;
end 13'h565:    begin Red = 8'h9a;    Green = 8'ha0;    Blue = 8'h96;
end 13'h566:    begin Red = 8'h78;    Green = 8'h8c;    Blue = 8'h7a;
end 13'h567:    begin Red = 8'h93;    Green = 8'h8e;    Blue = 8'h90;
end 13'h568:    begin Red = 8'h66;    Green = 8'h7a;    Blue = 8'h62;
end 13'h569:    begin Red = 8'h91;    Green = 8'h95;    Blue = 8'h92;
end 13'h56a:    begin Red = 8'h69;    Green = 8'h7d;    Blue = 8'h66;
end 13'h56b:    begin Red = 8'h71;    Green = 8'h79;    Blue = 8'h6c;
end 13'h56c:    begin Red = 8'h90;    Green = 8'h91;    Blue = 8'h8c;
end 13'h56d:    begin Red = 8'h94;    Green = 8'h92;    Blue = 8'h8c;
end 13'h56e:    begin Red = 8'hb1;    Green = 8'h98;    Blue = 8'h77;
end 13'h56f:    begin Red = 8'he1;    Green = 8'hc0;    Blue = 8'h9b;
end 13'h570:    begin Red = 8'hde;    Green = 8'hbf;    Blue = 8'h9f;
end 13'h571:    begin Red = 8'hdd;    Green = 8'hb3;    Blue = 8'h8b;
end 13'h572:    begin Red = 8'hd7;    Green = 8'hb0;    Blue = 8'h8e;
end 13'h573:    begin Red = 8'hd4;    Green = 8'hb4;    Blue = 8'h8b;
end 13'h574:    begin Red = 8'hd8;    Green = 8'hb3;    Blue = 8'h8c;
end 13'h575:    begin Red = 8'hd8;    Green = 8'haf;    Blue = 8'h89;
end 13'h576:    begin Red = 8'h9f;    Green = 8'h74;    Blue = 8'h55;
end 13'h577:    begin Red = 8'ha1;    Green = 8'h84;    Blue = 8'h5e;
end 13'h578:    begin Red = 8'h91;    Green = 8'h97;    Blue = 8'h7e;
end 13'h579:    begin Red = 8'h8e;    Green = 8'h8b;    Blue = 8'h88;
end 13'h57a:    begin Red = 8'hdb;    Green = 8'hb4;    Blue = 8'h88;
end 13'h57b:    begin Red = 8'h76;    Green = 8'h71;    Blue = 8'h5c;
end 13'h57c:    begin Red = 8'ha5;    Green = 8'hb7;    Blue = 8'h46;
end 13'h57d:    begin Red = 8'h7e;    Green = 8'h87;    Blue = 8'h65;
end 13'h57e:    begin Red = 8'hb7;    Green = 8'hd0;    Blue = 8'h46;
end 13'h57f:    begin Red = 8'hb0;    Green = 8'hc7;    Blue = 8'h51;
end 13'h580:    begin Red = 8'h3d;    Green = 8'h40;    Blue = 8'h3f;
end 13'h581:    begin Red = 8'h4f;    Green = 8'h56;    Blue = 8'h3f;
end 13'h582:    begin Red = 8'h54;    Green = 8'h70;    Blue = 8'h3a;
end 13'h583:    begin Red = 8'h5d;    Green = 8'h67;    Blue = 8'h3c;
end 13'h584:    begin Red = 8'h56;    Green = 8'h61;    Blue = 8'h39;
end 13'h585:    begin Red = 8'hb3;    Green = 8'ha6;    Blue = 8'h8b;
end 13'h586:    begin Red = 8'hb1;    Green = 8'h9a;    Blue = 8'h80;
end 13'h587:    begin Red = 8'hc9;    Green = 8'hb6;    Blue = 8'h93;
end 13'h588:    begin Red = 8'hdd;    Green = 8'hc1;    Blue = 8'ha1;
end 13'h589:    begin Red = 8'hcc;    Green = 8'haf;    Blue = 8'ha0;
end 13'h58a:    begin Red = 8'h56;    Green = 8'h61;    Blue = 8'h46;
end 13'h58b:    begin Red = 8'h53;    Green = 8'h57;    Blue = 8'h47;
end 13'h58c:    begin Red = 8'h52;    Green = 8'h5b;    Blue = 8'h43;
end 13'h58d:    begin Red = 8'h5e;    Green = 8'h68;    Blue = 8'h43;
end 13'h58e:    begin Red = 8'h85;    Green = 8'h7a;    Blue = 8'h63;
end 13'h58f:    begin Red = 8'h7b;    Green = 8'h78;    Blue = 8'h54;
end 13'h590:    begin Red = 8'h7e;    Green = 8'h7d;    Blue = 8'h5e;
end 13'h591:    begin Red = 8'heb;    Green = 8'hd3;    Blue = 8'hb5;
end 13'h592:    begin Red = 8'hdf;    Green = 8'hca;    Blue = 8'hb7;
end 13'h593:    begin Red = 8'he1;    Green = 8'hcd;    Blue = 8'had;
end 13'h594:    begin Red = 8'hed;    Green = 8'hd2;    Blue = 8'hb0;
end 13'h595:    begin Red = 8'hbf;    Green = 8'haf;    Blue = 8'h8c;
end 13'h596:    begin Red = 8'hde;    Green = 8'hcd;    Blue = 8'ha6;
end 13'h597:    begin Red = 8'he5;    Green = 8'hc6;    Blue = 8'ha7;
end 13'h598:    begin Red = 8'h98;    Green = 8'h97;    Blue = 8'h9b;
end 13'h599:    begin Red = 8'h95;    Green = 8'h9e;    Blue = 8'h99;
end 13'h59a:    begin Red = 8'h9b;    Green = 8'h9e;    Blue = 8'ha0;
end 13'h59b:    begin Red = 8'h9e;    Green = 8'h99;    Blue = 8'h9b;
end 13'h59c:    begin Red = 8'h7a;    Green = 8'h95;    Blue = 8'h7b;
end 13'h59d:    begin Red = 8'h97;    Green = 8'h9f;    Blue = 8'h9e;
end 13'h59e:    begin Red = 8'h72;    Green = 8'h7c;    Blue = 8'h6a;
end 13'h59f:    begin Red = 8'h65;    Green = 8'h7b;    Blue = 8'h5f;
end 13'h5a0:    begin Red = 8'h85;    Green = 8'h9c;    Blue = 8'h86;
end 13'h5a1:    begin Red = 8'h6e;    Green = 8'h7a;    Blue = 8'h69;
end 13'h5a2:    begin Red = 8'hac;    Green = 8'ha3;    Blue = 8'ha4;
end 13'h5a3:    begin Red = 8'h75;    Green = 8'h82;    Blue = 8'h6c;
end 13'h5a4:    begin Red = 8'h77;    Green = 8'h94;    Blue = 8'h86;
end 13'h5a5:    begin Red = 8'hb3;    Green = 8'h94;    Blue = 8'h75;
end 13'h5a6:    begin Red = 8'he2;    Green = 8'hc2;    Blue = 8'h9f;
end 13'h5a7:    begin Red = 8'h97;    Green = 8'h7b;    Blue = 8'h50;
end 13'h5a8:    begin Red = 8'ha0;    Green = 8'h79;    Blue = 8'h57;
end 13'h5a9:    begin Red = 8'hec;    Green = 8'hbe;    Blue = 8'h96;
end 13'h5aa:    begin Red = 8'he2;    Green = 8'hbe;    Blue = 8'h90;
end 13'h5ab:    begin Red = 8'he9;    Green = 8'hb9;    Blue = 8'h8e;
end 13'h5ac:    begin Red = 8'he9;    Green = 8'hbc;    Blue = 8'h8c;
end 13'h5ad:    begin Red = 8'he7;    Green = 8'hc0;    Blue = 8'h8c;
end 13'h5ae:    begin Red = 8'hf4;    Green = 8'hc4;    Blue = 8'h9b;
end 13'h5af:    begin Red = 8'h64;    Green = 8'h61;    Blue = 8'h42;
end 13'h5b0:    begin Red = 8'h7a;    Green = 8'h7a;    Blue = 8'h5d;
end 13'h5b1:    begin Red = 8'h80;    Green = 8'h7d;    Blue = 8'h66;
end 13'h5b2:    begin Red = 8'h83;    Green = 8'h79;    Blue = 8'h5a;
end 13'h5b3:    begin Red = 8'h5c;    Green = 8'h6e;    Blue = 8'h4b;
end 13'h5b4:    begin Red = 8'he1;    Green = 8'hb3;    Blue = 8'h8e;
end 13'h5b5:    begin Red = 8'hdb;    Green = 8'hb1;    Blue = 8'h8e;
end 13'h5b6:    begin Red = 8'h87;    Green = 8'h80;    Blue = 8'h5d;
end 13'h5b7:    begin Red = 8'h9f;    Green = 8'hac;    Blue = 8'h49;
end 13'h5b8:    begin Red = 8'h9b;    Green = 8'hab;    Blue = 8'h4f;
end 13'h5b9:    begin Red = 8'h88;    Green = 8'h97;    Blue = 8'h50;
end 13'h5ba:    begin Red = 8'h9b;    Green = 8'haf;    Blue = 8'h4e;
end 13'h5bb:    begin Red = 8'ha7;    Green = 8'hbe;    Blue = 8'h45;
end 13'h5bc:    begin Red = 8'h79;    Green = 8'h83;    Blue = 8'h5d;
end 13'h5bd:    begin Red = 8'had;    Green = 8'hc3;    Blue = 8'h54;
end 13'h5be:    begin Red = 8'h4a;    Green = 8'h4e;    Blue = 8'h45;
end 13'h5bf:    begin Red = 8'h60;    Green = 8'h68;    Blue = 8'h40;
end 13'h5c0:    begin Red = 8'h69;    Green = 8'h70;    Blue = 8'h42;
end 13'h5c1:    begin Red = 8'hb7;    Green = 8'h9a;    Blue = 8'h83;
end 13'h5c2:    begin Red = 8'hcd;    Green = 8'hba;    Blue = 8'h94;
end 13'h5c3:    begin Red = 8'hd9;    Green = 8'hbd;    Blue = 8'ha2;
end 13'h5c4:    begin Red = 8'h80;    Green = 8'h71;    Blue = 8'h5d;
end 13'h5c5:    begin Red = 8'hb8;    Green = 8'hac;    Blue = 8'h8d;
end 13'h5c6:    begin Red = 8'hbb;    Green = 8'hac;    Blue = 8'h90;
end 13'h5c7:    begin Red = 8'hbc;    Green = 8'haa;    Blue = 8'h88;
end 13'h5c8:    begin Red = 8'hb7;    Green = 8'ha4;    Blue = 8'h90;
end 13'h5c9:    begin Red = 8'hb6;    Green = 8'haa;    Blue = 8'h90;
end 13'h5ca:    begin Red = 8'hbb;    Green = 8'ha9;    Blue = 8'h96;
end 13'h5cb:    begin Red = 8'h60;    Green = 8'h62;    Blue = 8'h4a;
end 13'h5cc:    begin Red = 8'hd2;    Green = 8'hb3;    Blue = 8'h94;
end 13'h5cd:    begin Red = 8'he2;    Green = 8'hc7;    Blue = 8'had;
end 13'h5ce:    begin Red = 8'hdb;    Green = 8'hc7;    Blue = 8'haf;
end 13'h5cf:    begin Red = 8'ha0;    Green = 8'hb8;    Blue = 8'ha2;
end 13'h5d0:    begin Red = 8'h9a;    Green = 8'h95;    Blue = 8'h9d;
end 13'h5d1:    begin Red = 8'h95;    Green = 8'h9a;    Blue = 8'h97;
end 13'h5d2:    begin Red = 8'h7e;    Green = 8'h93;    Blue = 8'h75;
end 13'h5d3:    begin Red = 8'h9d;    Green = 8'h9c;    Blue = 8'h99;
end 13'h5d4:    begin Red = 8'h78;    Green = 8'h94;    Blue = 8'h79;
end 13'h5d5:    begin Red = 8'h98;    Green = 8'h7a;    Blue = 8'h59;
end 13'h5d6:    begin Red = 8'h98;    Green = 8'h7f;    Blue = 8'h58;
end 13'h5d7:    begin Red = 8'hd1;    Green = 8'hb7;    Blue = 8'h8c;
end 13'h5d8:    begin Red = 8'hd0;    Green = 8'hb7;    Blue = 8'h88;
end 13'h5d9:    begin Red = 8'h5a;    Green = 8'h67;    Blue = 8'h3e;
end 13'h5da:    begin Red = 8'h86;    Green = 8'h94;    Blue = 8'h65;
end 13'h5db:    begin Red = 8'h84;    Green = 8'h7e;    Blue = 8'h5f;
end 13'h5dc:    begin Red = 8'h7c;    Green = 8'h80;    Blue = 8'h5d;
end 13'h5dd:    begin Red = 8'h67;    Green = 8'h75;    Blue = 8'h53;
end 13'h5de:    begin Red = 8'hdc;    Green = 8'haf;    Blue = 8'h92;
end 13'h5df:    begin Red = 8'h7b;    Green = 8'h70;    Blue = 8'h5b;
end 13'h5e0:    begin Red = 8'h6b;    Green = 8'h66;    Blue = 8'h55;
end 13'h5e1:    begin Red = 8'h71;    Green = 8'h63;    Blue = 8'h53;
end 13'h5e2:    begin Red = 8'hb2;    Green = 8'hca;    Blue = 8'h40;
end 13'h5e3:    begin Red = 8'h7b;    Green = 8'h87;    Blue = 8'h53;
end 13'h5e4:    begin Red = 8'had;    Green = 8'hc1;    Blue = 8'h46;
end 13'h5e5:    begin Red = 8'hb3;    Green = 8'hcc;    Blue = 8'h4c;
end 13'h5e6:    begin Red = 8'haf;    Green = 8'hc7;    Blue = 8'h45;
end 13'h5e7:    begin Red = 8'h65;    Green = 8'h61;    Blue = 8'h4a;
end 13'h5e8:    begin Red = 8'hb9;    Green = 8'ha1;    Blue = 8'h8e;
end 13'h5e9:    begin Red = 8'h98;    Green = 8'h8a;    Blue = 8'h6d;
end 13'h5ea:    begin Red = 8'hfa;    Green = 8'he4;    Blue = 8'hc5;
end 13'h5eb:    begin Red = 8'hd9;    Green = 8'hc2;    Blue = 8'ha2;
end 13'h5ec:    begin Red = 8'h96;    Green = 8'h87;    Blue = 8'h6f;
end 13'h5ed:    begin Red = 8'h8e;    Green = 8'h78;    Blue = 8'h67;
end 13'h5ee:    begin Red = 8'h85;    Green = 8'h78;    Blue = 8'h69;
end 13'h5ef:    begin Red = 8'h8f;    Green = 8'h79;    Blue = 8'h6c;
end 13'h5f0:    begin Red = 8'ha7;    Green = 8'ha0;    Blue = 8'h57;
end 13'h5f1:    begin Red = 8'h6f;    Green = 8'h6e;    Blue = 8'h60;
end 13'h5f2:    begin Red = 8'had;    Green = 8'ha7;    Blue = 8'h4b;
end 13'h5f3:    begin Red = 8'ha4;    Green = 8'h9d;    Blue = 8'h53;
end 13'h5f4:    begin Red = 8'ha9;    Green = 8'ha8;    Blue = 8'h4c;
end 13'h5f5:    begin Red = 8'h9d;    Green = 8'h88;    Blue = 8'h6e;
end 13'h5f6:    begin Red = 8'ha7;    Green = 8'h98;    Blue = 8'h7d;
end 13'h5f7:    begin Red = 8'hb7;    Green = 8'ha1;    Blue = 8'h84;
end 13'h5f8:    begin Red = 8'h93;    Green = 8'hbd;    Blue = 8'h9a;
end 13'h5f9:    begin Red = 8'h9f;    Green = 8'hb5;    Blue = 8'h97;
end 13'h5fa:    begin Red = 8'h9b;    Green = 8'h97;    Blue = 8'ha0;
end 13'h5fb:    begin Red = 8'h7f;    Green = 8'h98;    Blue = 8'h8b;
end 13'h5fc:    begin Red = 8'h93;    Green = 8'ha8;    Blue = 8'h5b;
end 13'h5fd:    begin Red = 8'h98;    Green = 8'h9c;    Blue = 8'h3f;
end 13'h5fe:    begin Red = 8'ha4;    Green = 8'ha3;    Blue = 8'h4e;
end 13'h5ff:    begin Red = 8'ha3;    Green = 8'ha6;    Blue = 8'h54;
end 13'h600:    begin Red = 8'h83;    Green = 8'hb1;    Blue = 8'h82;
end 13'h601:    begin Red = 8'h88;    Green = 8'hb3;    Blue = 8'h7d;
end 13'h602:    begin Red = 8'h8a;    Green = 8'haf;    Blue = 8'h86;
end 13'h603:    begin Red = 8'h88;    Green = 8'hb0;    Blue = 8'h81;
end 13'h604:    begin Red = 8'h88;    Green = 8'h9b;    Blue = 8'h53;
end 13'h605:    begin Red = 8'h69;    Green = 8'h70;    Blue = 8'h5d;
end 13'h606:    begin Red = 8'ha6;    Green = 8'ha0;    Blue = 8'h4b;
end 13'h607:    begin Red = 8'h69;    Green = 8'h66;    Blue = 8'h52;
end 13'h608:    begin Red = 8'h69;    Green = 8'h5c;    Blue = 8'h54;
end 13'h609:    begin Red = 8'h5e;    Green = 8'h52;    Blue = 8'h56;
end 13'h60a:    begin Red = 8'h6c;    Green = 8'h69;    Blue = 8'h51;
end 13'h60b:    begin Red = 8'hb7;    Green = 8'hd0;    Blue = 8'h4e;
end 13'h60c:    begin Red = 8'h95;    Green = 8'ha9;    Blue = 8'h4b;
end 13'h60d:    begin Red = 8'ha7;    Green = 8'hbe;    Blue = 8'h4a;
end 13'h60e:    begin Red = 8'h67;    Green = 8'h53;    Blue = 8'h55;
end 13'h60f:    begin Red = 8'haa;    Green = 8'hc4;    Blue = 8'h3e;
end 13'h610:    begin Red = 8'h61;    Green = 8'h54;    Blue = 8'h59;
end 13'h611:    begin Red = 8'h94;    Green = 8'h89;    Blue = 8'h62;
end 13'h612:    begin Red = 8'h55;    Green = 8'h5a;    Blue = 8'h42;
end 13'h613:    begin Red = 8'h7d;    Green = 8'h8d;    Blue = 8'h45;
end 13'h614:    begin Red = 8'h6b;    Green = 8'h90;    Blue = 8'h48;
end 13'h615:    begin Red = 8'hd1;    Green = 8'hb7;    Blue = 8'h93;
end 13'h616:    begin Red = 8'ha1;    Green = 8'ha3;    Blue = 8'h41;
end 13'h617:    begin Red = 8'haa;    Green = 8'ha6;    Blue = 8'h48;
end 13'h618:    begin Red = 8'h83;    Green = 8'h80;    Blue = 8'h56;
end 13'h619:    begin Red = 8'hbd;    Green = 8'hde;    Blue = 8'h44;
end 13'h61a:    begin Red = 8'hb3;    Green = 8'hd6;    Blue = 8'h44;
end 13'h61b:    begin Red = 8'h9e;    Green = 8'hd2;    Blue = 8'h3c;
end 13'h61c:    begin Red = 8'hae;    Green = 8'hd5;    Blue = 8'h34;
end 13'h61d:    begin Red = 8'h90;    Green = 8'ha0;    Blue = 8'h4e;
end 13'h61e:    begin Red = 8'h8b;    Green = 8'h99;    Blue = 8'h56;
end 13'h61f:    begin Red = 8'h8e;    Green = 8'ha3;    Blue = 8'h52;
end 13'h620:    begin Red = 8'ha0;    Green = 8'hb7;    Blue = 8'h4e;
end 13'h621:    begin Red = 8'ha1;    Green = 8'hbe;    Blue = 8'h3d;
end 13'h622:    begin Red = 8'h79;    Green = 8'h78;    Blue = 8'h5a;
end 13'h623:    begin Red = 8'ha7;    Green = 8'haa;    Blue = 8'h4d;
end 13'h624:    begin Red = 8'hd1;    Green = 8'hca;    Blue = 8'h59;
end 13'h625:    begin Red = 8'h9b;    Green = 8'h9a;    Blue = 8'h48;
end 13'h626:    begin Red = 8'ha0;    Green = 8'h9d;    Blue = 8'h46;
end 13'h627:    begin Red = 8'ha0;    Green = 8'h8c;    Blue = 8'h6e;
end 13'h628:    begin Red = 8'hc7;    Green = 8'hc6;    Blue = 8'hd7;
end 13'h629:    begin Red = 8'hbe;    Green = 8'hb8;    Blue = 8'hc3;
end 13'h62a:    begin Red = 8'h9f;    Green = 8'hbc;    Blue = 8'h99;
end 13'h62b:    begin Red = 8'h9a;    Green = 8'hbe;    Blue = 8'h9d;
end 13'h62c:    begin Red = 8'h9c;    Green = 8'hbe;    Blue = 8'ha1;
end 13'h62d:    begin Red = 8'h88;    Green = 8'h90;    Blue = 8'h4b;
end 13'h62e:    begin Red = 8'h87;    Green = 8'h94;    Blue = 8'h48;
end 13'h62f:    begin Red = 8'h67;    Green = 8'h71;    Blue = 8'h34;
end 13'h630:    begin Red = 8'h72;    Green = 8'h76;    Blue = 8'h41;
end 13'h631:    begin Red = 8'h8c;    Green = 8'h90;    Blue = 8'h52;
end 13'h632:    begin Red = 8'h88;    Green = 8'h93;    Blue = 8'h4d;
end 13'h633:    begin Red = 8'ha0;    Green = 8'haf;    Blue = 8'h55;
end 13'h634:    begin Red = 8'h8c;    Green = 8'h96;    Blue = 8'h51;
end 13'h635:    begin Red = 8'h70;    Green = 8'h77;    Blue = 8'h43;
end 13'h636:    begin Red = 8'h9e;    Green = 8'hb0;    Blue = 8'h5a;
end 13'h637:    begin Red = 8'h95;    Green = 8'hac;    Blue = 8'h50;
end 13'h638:    begin Red = 8'h91;    Green = 8'hac;    Blue = 8'h53;
end 13'h639:    begin Red = 8'hce;    Green = 8'hb1;    Blue = 8'h8e;
end 13'h63a:    begin Red = 8'hc7;    Green = 8'ha3;    Blue = 8'h7d;
end 13'h63b:    begin Red = 8'hc3;    Green = 8'ha0;    Blue = 8'h84;
end 13'h63c:    begin Red = 8'h94;    Green = 8'ha0;    Blue = 8'h42;
end 13'h63d:    begin Red = 8'h9a;    Green = 8'ha2;    Blue = 8'h49;
end 13'h63e:    begin Red = 8'h75;    Green = 8'h7b;    Blue = 8'h61;
end 13'h63f:    begin Red = 8'h83;    Green = 8'h75;    Blue = 8'h51;
end 13'h640:    begin Red = 8'h73;    Green = 8'h6b;    Blue = 8'h57;
end 13'h641:    begin Red = 8'hb7;    Green = 8'hca;    Blue = 8'h3f;
end 13'h642:    begin Red = 8'h65;    Green = 8'h64;    Blue = 8'h61;
end 13'h643:    begin Red = 8'h78;    Green = 8'h77;    Blue = 8'h61;
end 13'h644:    begin Red = 8'ha4;    Green = 8'ha1;    Blue = 8'h54;
end 13'h645:    begin Red = 8'h6d;    Green = 8'h61;    Blue = 8'h4c;
end 13'h646:    begin Red = 8'h70;    Green = 8'h6a;    Blue = 8'h54;
end 13'h647:    begin Red = 8'h67;    Green = 8'h66;    Blue = 8'h4e;
end 13'h648:    begin Red = 8'ha7;    Green = 8'hc3;    Blue = 8'h4a;
end 13'h649:    begin Red = 8'h70;    Green = 8'h69;    Blue = 8'h59;
end 13'h64a:    begin Red = 8'h71;    Green = 8'h69;    Blue = 8'h4d;
end 13'h64b:    begin Red = 8'h8b;    Green = 8'h7d;    Blue = 8'h59;
end 13'h64c:    begin Red = 8'h59;    Green = 8'h65;    Blue = 8'h42;
end 13'h64d:    begin Red = 8'hb7;    Green = 8'ha0;    Blue = 8'h8c;
end 13'h64e:    begin Red = 8'hb1;    Green = 8'h9d;    Blue = 8'h84;
end 13'h64f:    begin Red = 8'h9a;    Green = 8'h85;    Blue = 8'h70;
end 13'h650:    begin Red = 8'hca;    Green = 8'hb0;    Blue = 8'h98;
end 13'h651:    begin Red = 8'h96;    Green = 8'h99;    Blue = 8'h3f;
end 13'h652:    begin Red = 8'h85;    Green = 8'h84;    Blue = 8'h5d;
end 13'h653:    begin Red = 8'h85;    Green = 8'h83;    Blue = 8'h61;
end 13'h654:    begin Red = 8'h87;    Green = 8'h7e;    Blue = 8'h5a;
end 13'h655:    begin Red = 8'hb4;    Green = 8'hd2;    Blue = 8'h47;
end 13'h656:    begin Red = 8'h86;    Green = 8'h97;    Blue = 8'h4d;
end 13'h657:    begin Red = 8'h6d;    Green = 8'h67;    Blue = 8'h5d;
end 13'h658:    begin Red = 8'h9d;    Green = 8'hb0;    Blue = 8'h41;
end 13'h659:    begin Red = 8'h80;    Green = 8'h7b;    Blue = 8'h56;
end 13'h65a:    begin Red = 8'hac;    Green = 8'ha3;    Blue = 8'h56;
end 13'h65b:    begin Red = 8'h9d;    Green = 8'h9a;    Blue = 8'h53;
end 13'h65c:    begin Red = 8'hca;    Green = 8'hc0;    Blue = 8'h61;
end 13'h65d:    begin Red = 8'h9f;    Green = 8'h89;    Blue = 8'h7a;
end 13'h65e:    begin Red = 8'h9e;    Green = 8'h8b;    Blue = 8'h6c;
end 13'h65f:    begin Red = 8'h98;    Green = 8'h83;    Blue = 8'h74;
end 13'h660:    begin Red = 8'hb1;    Green = 8'ha3;    Blue = 8'h81;
end 13'h661:    begin Red = 8'hbf;    Green = 8'hc2;    Blue = 8'hc9;
end 13'h662:    begin Red = 8'hbe;    Green = 8'hbe;    Blue = 8'hbe;
end 13'h663:    begin Red = 8'h72;    Green = 8'h70;    Blue = 8'h44;
end 13'h664:    begin Red = 8'h80;    Green = 8'h99;    Blue = 8'h88;
end 13'h665:    begin Red = 8'h8c;    Green = 8'h8e;    Blue = 8'h5a;
end 13'h666:    begin Red = 8'h9e;    Green = 8'hac;    Blue = 8'h5d;
end 13'h667:    begin Red = 8'h82;    Green = 8'h8c;    Blue = 8'h53;
end 13'h668:    begin Red = 8'h98;    Green = 8'hb3;    Blue = 8'h55;
end 13'h669:    begin Red = 8'hd4;    Green = 8'hb5;    Blue = 8'h96;
end 13'h66a:    begin Red = 8'hc9;    Green = 8'ha7;    Blue = 8'h80;
end 13'h66b:    begin Red = 8'hc9;    Green = 8'hab;    Blue = 8'h84;
end 13'h66c:    begin Red = 8'h9a;    Green = 8'ha1;    Blue = 8'h44;
end 13'h66d:    begin Red = 8'ha6;    Green = 8'ha3;    Blue = 8'h55;
end 13'h66e:    begin Red = 8'h7b;    Green = 8'h80;    Blue = 8'h58;
end 13'h66f:    begin Red = 8'h77;    Green = 8'h70;    Blue = 8'h62;
end 13'h670:    begin Red = 8'haa;    Green = 8'hc6;    Blue = 8'h4a;
end 13'h671:    begin Red = 8'hac;    Green = 8'hc1;    Blue = 8'h57;
end 13'h672:    begin Red = 8'hae;    Green = 8'hc1;    Blue = 8'h4b;
end 13'h673:    begin Red = 8'h8b;    Green = 8'h94;    Blue = 8'h57;
end 13'h674:    begin Red = 8'h89;    Green = 8'h84;    Blue = 8'h5f;
end 13'h675:    begin Red = 8'ha9;    Green = 8'ha0;    Blue = 8'h5b;
end 13'h676:    begin Red = 8'h71;    Green = 8'h6c;    Blue = 8'h52;
end 13'h677:    begin Red = 8'h6e;    Green = 8'h68;    Blue = 8'h57;
end 13'h678:    begin Red = 8'h63;    Green = 8'h5b;    Blue = 8'h51;
end 13'h679:    begin Red = 8'h65;    Green = 8'h5a;    Blue = 8'h55;
end 13'h67a:    begin Red = 8'h51;    Green = 8'h5f;    Blue = 8'h3e;
end 13'h67b:    begin Red = 8'hb3;    Green = 8'ha0;    Blue = 8'h7d;
end 13'h67c:    begin Red = 8'haf;    Green = 8'h9b;    Blue = 8'h7a;
end 13'h67d:    begin Red = 8'ha6;    Green = 8'h90;    Blue = 8'h72;
end 13'h67e:    begin Red = 8'hb1;    Green = 8'h9d;    Blue = 8'h7d;
end 13'h67f:    begin Red = 8'hd9;    Green = 8'hbb;    Blue = 8'ha9;
end 13'h680:    begin Red = 8'ha3;    Green = 8'ha2;    Blue = 8'h4b;
end 13'h681:    begin Red = 8'hb3;    Green = 8'hd6;    Blue = 8'h4a;
end 13'h682:    begin Red = 8'ha9;    Green = 8'hc5;    Blue = 8'h51;
end 13'h683:    begin Red = 8'hb8;    Green = 8'hd2;    Blue = 8'h48;
end 13'h684:    begin Red = 8'hab;    Green = 8'h94;    Blue = 8'h77;
end 13'h685:    begin Red = 8'hc4;    Green = 8'hbe;    Blue = 8'h55;
end 13'h686:    begin Red = 8'hc5;    Green = 8'hbe;    Blue = 8'h5a;
end 13'h687:    begin Red = 8'hc6;    Green = 8'hc3;    Blue = 8'h4a;
end 13'h688:    begin Red = 8'h9c;    Green = 8'h87;    Blue = 8'h71;
end 13'h689:    begin Red = 8'ha2;    Green = 8'ha6;    Blue = 8'hb5;
end 13'h68a:    begin Red = 8'ha7;    Green = 8'ha8;    Blue = 8'hac;
end 13'h68b:    begin Red = 8'hbb;    Green = 8'hbb;    Blue = 8'hbe;
end 13'h68c:    begin Red = 8'h88;    Green = 8'h9b;    Blue = 8'h99;
end 13'h68d:    begin Red = 8'h6e;    Green = 8'h80;    Blue = 8'h42;
end 13'h68e:    begin Red = 8'h79;    Green = 8'h95;    Blue = 8'h82;
end 13'h68f:    begin Red = 8'hb1;    Green = 8'h96;    Blue = 8'h7a;
end 13'h690:    begin Red = 8'he0;    Green = 8'hbc;    Blue = 8'h9b;
end 13'h691:    begin Red = 8'ha4;    Green = 8'ha8;    Blue = 8'h49;
end 13'h692:    begin Red = 8'h9f;    Green = 8'h9f;    Blue = 8'h51;
end 13'h693:    begin Red = 8'ha3;    Green = 8'ha0;    Blue = 8'h5a;
end 13'h694:    begin Red = 8'ha7;    Green = 8'ha3;    Blue = 8'h5a;
end 13'h695:    begin Red = 8'h7f;    Green = 8'h84;    Blue = 8'h5d;
end 13'h696:    begin Red = 8'h7a;    Green = 8'h6c;    Blue = 8'h5c;
end 13'h697:    begin Red = 8'hb2;    Green = 8'hca;    Blue = 8'h49;
end 13'h698:    begin Red = 8'h88;    Green = 8'h9b;    Blue = 8'h5d;
end 13'h699:    begin Red = 8'h8c;    Green = 8'h9c;    Blue = 8'h51;
end 13'h69a:    begin Red = 8'h9a;    Green = 8'hae;    Blue = 8'h49;
end 13'h69b:    begin Red = 8'hea;    Green = 8'hc1;    Blue = 8'h93;
end 13'h69c:    begin Red = 8'h7d;    Green = 8'h7b;    Blue = 8'h5c;
end 13'h69d:    begin Red = 8'ha4;    Green = 8'h9d;    Blue = 8'h4d;
end 13'h69e:    begin Red = 8'h66;    Green = 8'h65;    Blue = 8'h54;
end 13'h69f:    begin Red = 8'hb7;    Green = 8'hd9;    Blue = 8'h50;
end 13'h6a0:    begin Red = 8'h61;    Green = 8'h59;    Blue = 8'h4f;
end 13'h6a1:    begin Red = 8'ha3;    Green = 8'hc1;    Blue = 8'h3d;
end 13'h6a2:    begin Red = 8'ha7;    Green = 8'hcb;    Blue = 8'h3e;
end 13'h6a3:    begin Red = 8'ha3;    Green = 8'hc3;    Blue = 8'h39;
end 13'h6a4:    begin Red = 8'h6d;    Green = 8'h63;    Blue = 8'h54;
end 13'h6a5:    begin Red = 8'hcc;    Green = 8'hb3;    Blue = 8'ha3;
end 13'h6a6:    begin Red = 8'h97;    Green = 8'h92;    Blue = 8'h3a;
end 13'h6a7:    begin Red = 8'h9e;    Green = 8'h9b;    Blue = 8'h4e;
end 13'h6a8:    begin Red = 8'ha1;    Green = 8'h9b;    Blue = 8'h54;
end 13'h6a9:    begin Red = 8'hbe;    Green = 8'he0;    Blue = 8'h3f;
end 13'h6aa:    begin Red = 8'hba;    Green = 8'hd3;    Blue = 8'h4a;
end 13'h6ab:    begin Red = 8'h6a;    Green = 8'h61;    Blue = 8'h66;
end 13'h6ac:    begin Red = 8'h8b;    Green = 8'h92;    Blue = 8'h50;
end 13'h6ad:    begin Red = 8'ha6;    Green = 8'hbe;    Blue = 8'h3d;
end 13'h6ae:    begin Red = 8'h7c;    Green = 8'h84;    Blue = 8'h66;
end 13'h6af:    begin Red = 8'h7b;    Green = 8'h84;    Blue = 8'h62;
end 13'h6b0:    begin Red = 8'hac;    Green = 8'h98;    Blue = 8'h6c;
end 13'h6b1:    begin Red = 8'ha6;    Green = 8'ha7;    Blue = 8'h41;
end 13'h6b2:    begin Red = 8'h9b;    Green = 8'ha3;    Blue = 8'h46;
end 13'h6b3:    begin Red = 8'hcf;    Green = 8'hc8;    Blue = 8'h58;
end 13'h6b4:    begin Red = 8'hca;    Green = 8'hc4;    Blue = 8'h5a;
end 13'h6b5:    begin Red = 8'hcc;    Green = 8'hcc;    Blue = 8'h4e;
end 13'h6b6:    begin Red = 8'hb6;    Green = 8'h9f;    Blue = 8'h94;
end 13'h6b7:    begin Red = 8'h89;    Green = 8'h75;    Blue = 8'h65;
end 13'h6b8:    begin Red = 8'hc8;    Green = 8'hb1;    Blue = 8'h91;
end 13'h6b9:    begin Red = 8'hb5;    Green = 8'hb6;    Blue = 8'hb9;
end 13'h6ba:    begin Red = 8'hb7;    Green = 8'hb8;    Blue = 8'hbb;
end 13'h6bb:    begin Red = 8'h6c;    Green = 8'h75;    Blue = 8'h51;
end 13'h6bc:    begin Red = 8'h8f;    Green = 8'h9b;    Blue = 8'h65;
end 13'h6bd:    begin Red = 8'h8e;    Green = 8'h99;    Blue = 8'h5d;
end 13'h6be:    begin Red = 8'h86;    Green = 8'h9e;    Blue = 8'h88;
end 13'h6bf:    begin Red = 8'h87;    Green = 8'h9b;    Blue = 8'h93;
end 13'h6c0:    begin Red = 8'h8a;    Green = 8'h9e;    Blue = 8'h8f;
end 13'h6c1:    begin Red = 8'h7d;    Green = 8'h94;    Blue = 8'h48;
end 13'h6c2:    begin Red = 8'h94;    Green = 8'h9a;    Blue = 8'h47;
end 13'h6c3:    begin Red = 8'ha4;    Green = 8'ha3;    Blue = 8'h5d;
end 13'h6c4:    begin Red = 8'ha9;    Green = 8'ha9;    Blue = 8'h50;
end 13'h6c5:    begin Red = 8'h7f;    Green = 8'h82;    Blue = 8'h5a;
end 13'h6c6:    begin Red = 8'haf;    Green = 8'hd6;    Blue = 8'h49;
end 13'h6c7:    begin Red = 8'h67;    Green = 8'h69;    Blue = 8'h62;
end 13'h6c8:    begin Red = 8'he6;    Green = 8'hb9;    Blue = 8'h95;
end 13'h6c9:    begin Red = 8'ha0;    Green = 8'ha0;    Blue = 8'h42;
end 13'h6ca:    begin Red = 8'h6a;    Green = 8'h61;    Blue = 8'h51;
end 13'h6cb:    begin Red = 8'h88;    Green = 8'h7d;    Blue = 8'h57;
end 13'h6cc:    begin Red = 8'h8b;    Green = 8'h86;    Blue = 8'h56;
end 13'h6cd:    begin Red = 8'h88;    Green = 8'h7f;    Blue = 8'h52;
end 13'h6ce:    begin Red = 8'h88;    Green = 8'h7d;    Blue = 8'h5e;
end 13'h6cf:    begin Red = 8'h6e;    Green = 8'h78;    Blue = 8'h53;
end 13'h6d0:    begin Red = 8'ha0;    Green = 8'h86;    Blue = 8'h74;
end 13'h6d1:    begin Red = 8'hb3;    Green = 8'h9f;    Blue = 8'h8c;
end 13'h6d2:    begin Red = 8'hc7;    Green = 8'hac;    Blue = 8'h95;
end 13'h6d3:    begin Red = 8'hb9;    Green = 8'hb6;    Blue = 8'h36;
end 13'h6d4:    begin Red = 8'hc9;    Green = 8'hc0;    Blue = 8'h5a;
end 13'h6d5:    begin Red = 8'ha7;    Green = 8'h9a;    Blue = 8'h71;
end 13'h6d6:    begin Red = 8'ha7;    Green = 8'h92;    Blue = 8'h75;
end 13'h6d7:    begin Red = 8'h9f;    Green = 8'ha7;    Blue = 8'h3f;
end 13'h6d8:    begin Red = 8'hc7;    Green = 8'hb1;    Blue = 8'h8d;
end 13'h6d9:    begin Red = 8'h69;    Green = 8'h72;    Blue = 8'h51;
end 13'h6da:    begin Red = 8'h80;    Green = 8'h92;    Blue = 8'h8d;
end 13'h6db:    begin Red = 8'hde;    Green = 8'haf;    Blue = 8'h87;
end 13'h6dc:    begin Red = 8'hb7;    Green = 8'hc2;    Blue = 8'h49;
end 13'h6dd:    begin Red = 8'hc3;    Green = 8'hbf;    Blue = 8'h58;
end 13'h6de:    begin Red = 8'h9e;    Green = 8'h98;    Blue = 8'h58;
end 13'h6df:    begin Red = 8'hd9;    Green = 8'hb3;    Blue = 8'h84;
end 13'h6e0:    begin Red = 8'h6c;    Green = 8'h5f;    Blue = 8'h4a;
end 13'h6e1:    begin Red = 8'h51;    Green = 8'h52;    Blue = 8'h3f;
end 13'h6e2:    begin Red = 8'h65;    Green = 8'h58;    Blue = 8'h3b;
end 13'h6e3:    begin Red = 8'h6c;    Green = 8'h5d;    Blue = 8'h46;
end 13'h6e4:    begin Red = 8'hb3;    Green = 8'h90;    Blue = 8'h71;
end 13'h6e5:    begin Red = 8'h64;    Green = 8'h5c;    Blue = 8'h40;
end 13'h6e6:    begin Red = 8'h5f;    Green = 8'h5b;    Blue = 8'h44;
end 13'h6e7:    begin Red = 8'h75;    Green = 8'h77;    Blue = 8'h50;
end 13'h6e8:    begin Red = 8'hea;    Green = 8'hd7;    Blue = 8'hb4;
end 13'h6e9:    begin Red = 8'hfe;    Green = 8'he6;    Blue = 8'hc8;
end 13'h6ea:    begin Red = 8'hce;    Green = 8'hcb;    Blue = 8'h55;
end 13'h6eb:    begin Red = 8'hc9;    Green = 8'hc2;    Blue = 8'h55;
end 13'h6ec:    begin Red = 8'h7d;    Green = 8'h88;    Blue = 8'h55;
end 13'h6ed:    begin Red = 8'ha0;    Green = 8'hb7;    Blue = 8'h3c;
end 13'h6ee:    begin Red = 8'h9e;    Green = 8'hb0;    Blue = 8'h53;
end 13'h6ef:    begin Red = 8'h4e;    Green = 8'h51;    Blue = 8'h46;
end 13'h6f0:    begin Red = 8'he8;    Green = 8'hd5;    Blue = 8'haf;
end 13'h6f1:    begin Red = 8'heb;    Green = 8'hd2;    Blue = 8'hbc;
end 13'h6f2:    begin Red = 8'ha5;    Green = 8'h96;    Blue = 8'h67;
end 13'h6f3:    begin Red = 8'hef;    Green = 8'hd6;    Blue = 8'hb3;
end 13'h6f4:    begin Red = 8'he6;    Green = 8'hd4;    Blue = 8'h9f;
end 13'h6f5:    begin Red = 8'h9a;    Green = 8'ha0;    Blue = 8'hab;
end 13'h6f6:    begin Red = 8'ha2;    Green = 8'ha6;    Blue = 8'ha8;
end 13'h6f7:    begin Red = 8'hb9;    Green = 8'hbd;    Blue = 8'hbf;
end 13'h6f8:    begin Red = 8'hbc;    Green = 8'hbd;    Blue = 8'hc1;
end 13'h6f9:    begin Red = 8'h5e;    Green = 8'h62;    Blue = 8'h5d;
end 13'h6fa:    begin Red = 8'h6c;    Green = 8'h70;    Blue = 8'h62;
end 13'h6fb:    begin Red = 8'ha0;    Green = 8'hb0;    Blue = 8'h46;
end 13'h6fc:    begin Red = 8'ha2;    Green = 8'ha0;    Blue = 8'h4e;
end 13'h6fd:    begin Red = 8'ha7;    Green = 8'ha3;    Blue = 8'h50;
end 13'h6fe:    begin Red = 8'h84;    Green = 8'h81;    Blue = 8'h63;
end 13'h6ff:    begin Red = 8'haf;    Green = 8'hbe;    Blue = 8'h50;
end 13'h700:    begin Red = 8'h5e;    Green = 8'h5d;    Blue = 8'h46;
end 13'h701:    begin Red = 8'h41;    Green = 8'h52;    Blue = 8'h34;
end 13'h702:    begin Red = 8'hd9;    Green = 8'hb7;    Blue = 8'h8e;
end 13'h703:    begin Red = 8'h53;    Green = 8'h55;    Blue = 8'h40;
end 13'h704:    begin Red = 8'hc8;    Green = 8'h9e;    Blue = 8'h73;
end 13'h705:    begin Red = 8'h4f;    Green = 8'h53;    Blue = 8'h3b;
end 13'h706:    begin Red = 8'h54;    Green = 8'h50;    Blue = 8'h40;
end 13'h707:    begin Red = 8'h89;    Green = 8'h81;    Blue = 8'h5a;
end 13'h708:    begin Red = 8'h76;    Green = 8'h77;    Blue = 8'h54;
end 13'h709:    begin Red = 8'hb9;    Green = 8'h9a;    Blue = 8'h6b;
end 13'h70a:    begin Red = 8'h6c;    Green = 8'h5f;    Blue = 8'h42;
end 13'h70b:    begin Red = 8'h4e;    Green = 8'h59;    Blue = 8'h36;
end 13'h70c:    begin Red = 8'h88;    Green = 8'h9f;    Blue = 8'h5b;
end 13'h70d:    begin Red = 8'h95;    Green = 8'h80;    Blue = 8'h65;
end 13'h70e:    begin Red = 8'hd6;    Green = 8'hc1;    Blue = 8'h9b;
end 13'h70f:    begin Red = 8'h9a;    Green = 8'h87;    Blue = 8'h74;
end 13'h710:    begin Red = 8'hd2;    Green = 8'hd1;    Blue = 8'h4a;
end 13'h711:    begin Red = 8'h9b;    Green = 8'h98;    Blue = 8'h61;
end 13'h712:    begin Red = 8'h81;    Green = 8'h87;    Blue = 8'h5c;
end 13'h713:    begin Red = 8'h7b;    Green = 8'h76;    Blue = 8'h5b;
end 13'h714:    begin Red = 8'hb0;    Green = 8'hc6;    Blue = 8'h55;
end 13'h715:    begin Red = 8'ha4;    Green = 8'hbb;    Blue = 8'h47;
end 13'h716:    begin Red = 8'hbc;    Green = 8'h9b;    Blue = 8'h88;
end 13'h717:    begin Red = 8'hb3;    Green = 8'h98;    Blue = 8'h7e;
end 13'h718:    begin Red = 8'hff;    Green = 8'he9;    Blue = 8'hc3;
end 13'h719:    begin Red = 8'hff;    Green = 8'he2;    Blue = 8'hbf;
end 13'h71a:    begin Red = 8'h95;    Green = 8'h9d;    Blue = 8'ha5;
end 13'h71b:    begin Red = 8'h9b;    Green = 8'ha5;    Blue = 8'ha3;
end 13'h71c:    begin Red = 8'hb7;    Green = 8'hc3;    Blue = 8'hc1;
end 13'h71d:    begin Red = 8'h92;    Green = 8'hae;    Blue = 8'h94;
end 13'h71e:    begin Red = 8'h81;    Green = 8'h99;    Blue = 8'h91;
end 13'h71f:    begin Red = 8'h79;    Green = 8'h80;    Blue = 8'h55;
end 13'h720:    begin Red = 8'ha0;    Green = 8'hb5;    Blue = 8'h5a;
end 13'h721:    begin Red = 8'h7f;    Green = 8'h8f;    Blue = 8'h90;
end 13'h722:    begin Red = 8'h75;    Green = 8'h92;    Blue = 8'h8a;
end 13'h723:    begin Red = 8'he3;    Green = 8'hbf;    Blue = 8'h9e;
end 13'h724:    begin Red = 8'hdd;    Green = 8'hb7;    Blue = 8'h90;
end 13'h725:    begin Red = 8'hc9;    Green = 8'hc6;    Blue = 8'h4f;
end 13'h726:    begin Red = 8'hcd;    Green = 8'hc3;    Blue = 8'h5d;
end 13'h727:    begin Red = 8'h9b;    Green = 8'h98;    Blue = 8'h5a;
end 13'h728:    begin Red = 8'hb4;    Green = 8'hcb;    Blue = 8'h51;
end 13'h729:    begin Red = 8'ha3;    Green = 8'hb7;    Blue = 8'h4c;
end 13'h72a:    begin Red = 8'h5b;    Green = 8'h65;    Blue = 8'h46;
end 13'h72b:    begin Red = 8'hec;    Green = 8'hbd;    Blue = 8'h9a;
end 13'h72c:    begin Red = 8'hf1;    Green = 8'hbe;    Blue = 8'h9a;
end 13'h72d:    begin Red = 8'h62;    Green = 8'h5c;    Blue = 8'h4b;
end 13'h72e:    begin Red = 8'h6b;    Green = 8'h5a;    Blue = 8'h42;
end 13'h72f:    begin Red = 8'hb1;    Green = 8'h8f;    Blue = 8'h66;
end 13'h730:    begin Red = 8'hc1;    Green = 8'h97;    Blue = 8'h75;
end 13'h731:    begin Red = 8'hb9;    Green = 8'h94;    Blue = 8'h69;
end 13'h732:    begin Red = 8'h85;    Green = 8'h7b;    Blue = 8'h58;
end 13'h733:    begin Red = 8'haf;    Green = 8'h95;    Blue = 8'h6e;
end 13'h734:    begin Red = 8'hb9;    Green = 8'h96;    Blue = 8'h6f;
end 13'h735:    begin Red = 8'hc4;    Green = 8'h91;    Blue = 8'h7b;
end 13'h736:    begin Red = 8'hb7;    Green = 8'h8e;    Blue = 8'h6f;
end 13'h737:    begin Red = 8'h68;    Green = 8'h63;    Blue = 8'h3d;
end 13'h738:    begin Red = 8'h63;    Green = 8'h5e;    Blue = 8'h43;
end 13'h739:    begin Red = 8'h65;    Green = 8'h5b;    Blue = 8'h46;
end 13'h73a:    begin Red = 8'h57;    Green = 8'h54;    Blue = 8'h3d;
end 13'h73b:    begin Red = 8'ha3;    Green = 8'h8e;    Blue = 8'h6c;
end 13'h73c:    begin Red = 8'h63;    Green = 8'h76;    Blue = 8'h46;
end 13'h73d:    begin Red = 8'h98;    Green = 8'h83;    Blue = 8'h67;
end 13'h73e:    begin Red = 8'hed;    Green = 8'hd8;    Blue = 8'hb1;
end 13'h73f:    begin Red = 8'hd9;    Green = 8'hc4;    Blue = 8'h9b;
end 13'h740:    begin Red = 8'h96;    Green = 8'h8b;    Blue = 8'h75;
end 13'h741:    begin Red = 8'ha1;    Green = 8'ha2;    Blue = 8'h58;
end 13'h742:    begin Red = 8'h9b;    Green = 8'hb2;    Blue = 8'h4c;
end 13'h743:    begin Red = 8'hab;    Green = 8'hc0;    Blue = 8'h51;
end 13'h744:    begin Red = 8'hb3;    Green = 8'hce;    Blue = 8'h42;
end 13'h745:    begin Red = 8'hc0;    Green = 8'hda;    Blue = 8'h4e;
end 13'h746:    begin Red = 8'hb5;    Green = 8'hbb;    Blue = 8'hc4;
end 13'h747:    begin Red = 8'hb7;    Green = 8'hc9;    Blue = 8'hbc;
end 13'h748:    begin Red = 8'hce;    Green = 8'h94;    Blue = 8'hc4;
end 13'h749:    begin Red = 8'hd1;    Green = 8'h96;    Blue = 8'hb3;
end 13'h74a:    begin Red = 8'hca;    Green = 8'h9a;    Blue = 8'hc3;
end 13'h74b:    begin Red = 8'hd5;    Green = 8'he1;    Blue = 8'hdb;
end 13'h74c:    begin Red = 8'hd9;    Green = 8'hcd;    Blue = 8'hb2;
end 13'h74d:    begin Red = 8'h89;    Green = 8'h9d;    Blue = 8'h55;
end 13'h74e:    begin Red = 8'h58;    Green = 8'h5e;    Blue = 8'h3f;
end 13'h74f:    begin Red = 8'h9b;    Green = 8'hb6;    Blue = 8'h3f;
end 13'h750:    begin Red = 8'hc5;    Green = 8'hac;    Blue = 8'h7e;
end 13'h751:    begin Red = 8'hab;    Green = 8'h9b;    Blue = 8'h55;
end 13'h752:    begin Red = 8'hca;    Green = 8'hc1;    Blue = 8'h5d;
end 13'h753:    begin Red = 8'ha0;    Green = 8'h9f;    Blue = 8'h55;
end 13'h754:    begin Red = 8'h7b;    Green = 8'h78;    Blue = 8'h64;
end 13'h755:    begin Red = 8'h80;    Green = 8'h84;    Blue = 8'h57;
end 13'h756:    begin Red = 8'h85;    Green = 8'h79;    Blue = 8'h4e;
end 13'h757:    begin Red = 8'h63;    Green = 8'h5d;    Blue = 8'h47;
end 13'h758:    begin Red = 8'h5b;    Green = 8'h55;    Blue = 8'h3f;
end 13'h759:    begin Red = 8'h57;    Green = 8'h55;    Blue = 8'h42;
end 13'h75a:    begin Red = 8'hbc;    Green = 8'h9d;    Blue = 8'h70;
end 13'h75b:    begin Red = 8'hd2;    Green = 8'h99;    Blue = 8'h78;
end 13'h75c:    begin Red = 8'h5e;    Green = 8'h55;    Blue = 8'h42;
end 13'h75d:    begin Red = 8'h83;    Green = 8'h78;    Blue = 8'h55;
end 13'h75e:    begin Red = 8'h62;    Green = 8'h51;    Blue = 8'h42;
end 13'h75f:    begin Red = 8'h54;    Green = 8'h57;    Blue = 8'h3d;
end 13'h760:    begin Red = 8'h69;    Green = 8'h5f;    Blue = 8'h4c;
end 13'h761:    begin Red = 8'h8b;    Green = 8'h7e;    Blue = 8'h4d;
end 13'h762:    begin Red = 8'h8b;    Green = 8'h7f;    Blue = 8'h48;
end 13'h763:    begin Red = 8'h8a;    Green = 8'h79;    Blue = 8'h47;
end 13'h764:    begin Red = 8'h81;    Green = 8'h78;    Blue = 8'h4e;
end 13'h765:    begin Red = 8'h73;    Green = 8'h72;    Blue = 8'h3f;
end 13'h766:    begin Red = 8'hff;    Green = 8'he2;    Blue = 8'hc5;
end 13'h767:    begin Red = 8'hbe;    Green = 8'ha3;    Blue = 8'h93;
end 13'h768:    begin Red = 8'h7d;    Green = 8'h68;    Blue = 8'h62;
end 13'h769:    begin Red = 8'hd9;    Green = 8'hc1;    Blue = 8'hab;
end 13'h76a:    begin Red = 8'h9b;    Green = 8'h86;    Blue = 8'h77;
end 13'h76b:    begin Red = 8'hdf;    Green = 8'hc5;    Blue = 8'hbf;
end 13'h76c:    begin Red = 8'hd8;    Green = 8'hb8;    Blue = 8'hc1;
end 13'h76d:    begin Red = 8'hce;    Green = 8'hc3;    Blue = 8'h61;
end 13'h76e:    begin Red = 8'h9b;    Green = 8'h94;    Blue = 8'h4b;
end 13'h76f:    begin Red = 8'hd6;    Green = 8'hca;    Blue = 8'h5e;
end 13'h770:    begin Red = 8'hb7;    Green = 8'had;    Blue = 8'h54;
end 13'h771:    begin Red = 8'h76;    Green = 8'h74;    Blue = 8'h5a;
end 13'h772:    begin Red = 8'hac;    Green = 8'hc9;    Blue = 8'h43;
end 13'h773:    begin Red = 8'h57;    Green = 8'h49;    Blue = 8'h5d;
end 13'h774:    begin Red = 8'hb5;    Green = 8'hcd;    Blue = 8'h4e;
end 13'h775:    begin Red = 8'h7d;    Green = 8'h87;    Blue = 8'h5a;
end 13'h776:    begin Red = 8'h46;    Green = 8'h4d;    Blue = 8'h3c;
end 13'h777:    begin Red = 8'h79;    Green = 8'h86;    Blue = 8'h4c;
end 13'h778:    begin Red = 8'hf9;    Green = 8'hd5;    Blue = 8'hb6;
end 13'h779:    begin Red = 8'hbe;    Green = 8'h78;    Blue = 8'haf;
end 13'h77a:    begin Red = 8'hb6;    Green = 8'h76;    Blue = 8'haf;
end 13'h77b:    begin Red = 8'hd2;    Green = 8'he4;    Blue = 8'hda;
end 13'h77c:    begin Red = 8'hd2;    Green = 8'he2;    Blue = 8'he7;
end 13'h77d:    begin Red = 8'hd2;    Green = 8'hd9;    Blue = 8'hd5;
end 13'h77e:    begin Red = 8'hd1;    Green = 8'hd3;    Blue = 8'hd7;
end 13'h77f:    begin Red = 8'hf4;    Green = 8'hed;    Blue = 8'hd2;
end 13'h780:    begin Red = 8'hf3;    Green = 8'hed;    Blue = 8'hca;
end 13'h781:    begin Red = 8'hd6;    Green = 8'hcf;    Blue = 8'had;
end 13'h782:    begin Red = 8'hd9;    Green = 8'hd8;    Blue = 8'had;
end 13'h783:    begin Red = 8'hab;    Green = 8'hc0;    Blue = 8'ha4;
end 13'h784:    begin Red = 8'h7d;    Green = 8'h9a;    Blue = 8'h84;
end 13'h785:    begin Red = 8'h88;    Green = 8'h9c;    Blue = 8'h8d;
end 13'h786:    begin Red = 8'h80;    Green = 8'h89;    Blue = 8'h58;
end 13'h787:    begin Red = 8'h6d;    Green = 8'h6e;    Blue = 8'h6a;
end 13'h788:    begin Red = 8'h8c;    Green = 8'ha3;    Blue = 8'h4f;
end 13'h789:    begin Red = 8'h84;    Green = 8'h95;    Blue = 8'h60;
end 13'h78a:    begin Red = 8'h85;    Green = 8'h92;    Blue = 8'h92;
end 13'h78b:    begin Red = 8'h7d;    Green = 8'h8f;    Blue = 8'h8d;
end 13'h78c:    begin Red = 8'h71;    Green = 8'h8d;    Blue = 8'h88;
end 13'h78d:    begin Red = 8'he4;    Green = 8'hb8;    Blue = 8'h98;
end 13'h78e:    begin Red = 8'he4;    Green = 8'hb4;    Blue = 8'h97;
end 13'h78f:    begin Red = 8'hd3;    Green = 8'hc1;    Blue = 8'h5b;
end 13'h790:    begin Red = 8'h9e;    Green = 8'h96;    Blue = 8'h4f;
end 13'h791:    begin Red = 8'h9b;    Green = 8'h9d;    Blue = 8'h4e;
end 13'h792:    begin Red = 8'ha2;    Green = 8'ha6;    Blue = 8'h5b;
end 13'h793:    begin Red = 8'ha6;    Green = 8'h9d;    Blue = 8'h5d;
end 13'h794:    begin Red = 8'h62;    Green = 8'h5d;    Blue = 8'h55;
end 13'h795:    begin Red = 8'h3e;    Green = 8'h40;    Blue = 8'h44;
end 13'h796:    begin Red = 8'h87;    Green = 8'h7a;    Blue = 8'h4b;
end 13'h797:    begin Red = 8'hb7;    Green = 8'h8c;    Blue = 8'h73;
end 13'h798:    begin Red = 8'hc6;    Green = 8'h9b;    Blue = 8'h7a;
end 13'h799:    begin Red = 8'h8f;    Green = 8'h88;    Blue = 8'h5c;
end 13'h79a:    begin Red = 8'h69;    Green = 8'h5e;    Blue = 8'h43;
end 13'h79b:    begin Red = 8'h8a;    Green = 8'h74;    Blue = 8'h4c;
end 13'h79c:    begin Red = 8'h82;    Green = 8'h75;    Blue = 8'h4c;
end 13'h79d:    begin Red = 8'hf1;    Green = 8'hd5;    Blue = 8'hbb;
end 13'h79e:    begin Red = 8'hc1;    Green = 8'ha1;    Blue = 8'h99;
end 13'h79f:    begin Red = 8'h98;    Green = 8'h8b;    Blue = 8'h78;
end 13'h7a0:    begin Red = 8'hd6;    Green = 8'hc1;    Blue = 8'ha7;
end 13'h7a1:    begin Red = 8'hce;    Green = 8'hb4;    Blue = 8'ha8;
end 13'h7a2:    begin Red = 8'hc6;    Green = 8'hbc;    Blue = 8'h5e;
end 13'h7a3:    begin Red = 8'hcf;    Green = 8'hc9;    Blue = 8'h5c;
end 13'h7a4:    begin Red = 8'hac;    Green = 8'hbe;    Blue = 8'h45;
end 13'h7a5:    begin Red = 8'h61;    Green = 8'h55;    Blue = 8'h55;
end 13'h7a6:    begin Red = 8'hb3;    Green = 8'hc1;    Blue = 8'h55;
end 13'h7a7:    begin Red = 8'h69;    Green = 8'h69;    Blue = 8'h4d;
end 13'h7a8:    begin Red = 8'h69;    Green = 8'h77;    Blue = 8'h51;
end 13'h7a9:    begin Red = 8'h90;    Green = 8'h94;    Blue = 8'h61;
end 13'h7aa:    begin Red = 8'hff;    Green = 8'hd4;    Blue = 8'hc1;
end 13'h7ab:    begin Red = 8'hbf;    Green = 8'h89;    Blue = 8'hb2;
end 13'h7ac:    begin Red = 8'hb3;    Green = 8'h76;    Blue = 8'hac;
end 13'h7ad:    begin Red = 8'hcc;    Green = 8'hd2;    Blue = 8'hd5;
end 13'h7ae:    begin Red = 8'hd6;    Green = 8'hd5;    Blue = 8'hd9;
end 13'h7af:    begin Red = 8'hed;    Green = 8'hea;    Blue = 8'hca;
end 13'h7b0:    begin Red = 8'h83;    Green = 8'h99;    Blue = 8'h8e;
end 13'h7b1:    begin Red = 8'hc4;    Green = 8'hbb;    Blue = 8'h59;
end 13'h7b2:    begin Red = 8'h9d;    Green = 8'ha0;    Blue = 8'h4c;
end 13'h7b3:    begin Red = 8'h9a;    Green = 8'h99;    Blue = 8'h4f;
end 13'h7b4:    begin Red = 8'hca;    Green = 8'hbe;    Blue = 8'h68;
end 13'h7b5:    begin Red = 8'haa;    Green = 8'ha7;    Blue = 8'h5a;
end 13'h7b6:    begin Red = 8'h87;    Green = 8'h7f;    Blue = 8'h62;
end 13'h7b7:    begin Red = 8'hbe;    Green = 8'hd6;    Blue = 8'h48;
end 13'h7b8:    begin Red = 8'h6d;    Green = 8'h6c;    Blue = 8'h4e;
end 13'h7b9:    begin Red = 8'h84;    Green = 8'h92;    Blue = 8'h4f;
end 13'h7ba:    begin Red = 8'haa;    Green = 8'hbc;    Blue = 8'h4a;
end 13'h7bb:    begin Red = 8'had;    Green = 8'hce;    Blue = 8'h39;
end 13'h7bc:    begin Red = 8'hae;    Green = 8'hc4;    Blue = 8'h43;
end 13'h7bd:    begin Red = 8'h4a;    Green = 8'h4d;    Blue = 8'h3e;
end 13'h7be:    begin Red = 8'h62;    Green = 8'h59;    Blue = 8'h47;
end 13'h7bf:    begin Red = 8'hc6;    Green = 8'h94;    Blue = 8'h71;
end 13'h7c0:    begin Red = 8'hb0;    Green = 8'h93;    Blue = 8'h69;
end 13'h7c1:    begin Red = 8'h86;    Green = 8'h75;    Blue = 8'h46;
end 13'h7c2:    begin Red = 8'h65;    Green = 8'h5b;    Blue = 8'h3d;
end 13'h7c3:    begin Red = 8'h88;    Green = 8'h7a;    Blue = 8'h4f;
end 13'h7c4:    begin Red = 8'h7e;    Green = 8'h71;    Blue = 8'h47;
end 13'h7c5:    begin Red = 8'he4;    Green = 8'hc9;    Blue = 8'hac;
end 13'h7c6:    begin Red = 8'hf3;    Green = 8'hd7;    Blue = 8'hb7;
end 13'h7c7:    begin Red = 8'h83;    Green = 8'h71;    Blue = 8'h64;
end 13'h7c8:    begin Red = 8'h89;    Green = 8'h7f;    Blue = 8'h65;
end 13'h7c9:    begin Red = 8'hf5;    Green = 8'he5;    Blue = 8'hbd;
end 13'h7ca:    begin Red = 8'h92;    Green = 8'h94;    Blue = 8'h3a;
end 13'h7cb:    begin Red = 8'hc5;    Green = 8'hc1;    Blue = 8'h5d;
end 13'h7cc:    begin Red = 8'h69;    Green = 8'h6c;    Blue = 8'h53;
end 13'h7cd:    begin Red = 8'h98;    Green = 8'hae;    Blue = 8'h3e;
end 13'h7ce:    begin Red = 8'h6e;    Green = 8'h66;    Blue = 8'h4a;
end 13'h7cf:    begin Red = 8'ha0;    Green = 8'hbe;    Blue = 8'h46;
end 13'h7d0:    begin Red = 8'h88;    Green = 8'h82;    Blue = 8'h57;
end 13'h7d1:    begin Red = 8'h61;    Green = 8'h68;    Blue = 8'h46;
end 13'h7d2:    begin Red = 8'hc1;    Green = 8'h8b;    Blue = 8'hb3;
end 13'h7d3:    begin Red = 8'hb7;    Green = 8'h7b;    Blue = 8'ha8;
end 13'h7d4:    begin Red = 8'hce;    Green = 8'hd9;    Blue = 8'hd3;
end 13'h7d5:    begin Red = 8'hcc;    Green = 8'h92;    Blue = 8'hbc;
end 13'h7d6:    begin Red = 8'hd1;    Green = 8'h9b;    Blue = 8'hc2;
end 13'h7d7:    begin Red = 8'he7;    Green = 8'he1;    Blue = 8'hc2;
end 13'h7d8:    begin Red = 8'hce;    Green = 8'hc7;    Blue = 8'ha8;
end 13'h7d9:    begin Red = 8'hd2;    Green = 8'hcd;    Blue = 8'haa;
end 13'h7da:    begin Red = 8'h54;    Green = 8'h5c;    Blue = 8'h34;
end 13'h7db:    begin Red = 8'h7b;    Green = 8'h7e;    Blue = 8'h61;
end 13'h7dc:    begin Red = 8'hd7;    Green = 8'hb5;    Blue = 8'h89;
end 13'h7dd:    begin Red = 8'h99;    Green = 8'h9b;    Blue = 8'h46;
end 13'h7de:    begin Red = 8'hc6;    Green = 8'hba;    Blue = 8'h5b;
end 13'h7df:    begin Red = 8'haa;    Green = 8'ha3;    Blue = 8'h52;
end 13'h7e0:    begin Red = 8'h84;    Green = 8'h84;    Blue = 8'h56;
end 13'h7e1:    begin Red = 8'h6c;    Green = 8'h65;    Blue = 8'h4f;
end 13'h7e2:    begin Red = 8'h71;    Green = 8'h67;    Blue = 8'h55;
end 13'h7e3:    begin Red = 8'hbb;    Green = 8'hd8;    Blue = 8'h4f;
end 13'h7e4:    begin Red = 8'h6b;    Green = 8'h68;    Blue = 8'h4a;
end 13'h7e5:    begin Red = 8'h8e;    Green = 8'h80;    Blue = 8'h55;
end 13'h7e6:    begin Red = 8'h63;    Green = 8'h65;    Blue = 8'h47;
end 13'h7e7:    begin Red = 8'hac;    Green = 8'h87;    Blue = 8'h58;
end 13'h7e8:    begin Red = 8'ha2;    Green = 8'h83;    Blue = 8'h54;
end 13'h7e9:    begin Red = 8'h5f;    Green = 8'h56;    Blue = 8'h3f;
end 13'h7ea:    begin Red = 8'h5a;    Green = 8'h5b;    Blue = 8'h40;
end 13'h7eb:    begin Red = 8'h84;    Green = 8'h72;    Blue = 8'h49;
end 13'h7ec:    begin Red = 8'ha1;    Green = 8'h79;    Blue = 8'h51;
end 13'h7ed:    begin Red = 8'h9e;    Green = 8'h78;    Blue = 8'h4f;
end 13'h7ee:    begin Red = 8'h9b;    Green = 8'h78;    Blue = 8'h4c;
end 13'h7ef:    begin Red = 8'h75;    Green = 8'h69;    Blue = 8'h5c;
end 13'h7f0:    begin Red = 8'h6e;    Green = 8'h5d;    Blue = 8'h4e;
end 13'h7f1:    begin Red = 8'hd6;    Green = 8'hd0;    Blue = 8'h59;
end 13'h7f2:    begin Red = 8'h5d;    Green = 8'h6c;    Blue = 8'h48;
end 13'h7f3:    begin Red = 8'hc0;    Green = 8'hbf;    Blue = 8'h5a;
end 13'h7f4:    begin Red = 8'hd9;    Green = 8'hcd;    Blue = 8'h60;
end 13'h7f5:    begin Red = 8'he7;    Green = 8'hdb;    Blue = 8'h5a;
end 13'h7f6:    begin Red = 8'h5d;    Green = 8'h48;    Blue = 8'h5f;
end 13'h7f7:    begin Red = 8'h67;    Green = 8'h58;    Blue = 8'h53;
end 13'h7f8:    begin Red = 8'ha2;    Green = 8'hbc;    Blue = 8'h4a;
end 13'h7f9:    begin Red = 8'hac;    Green = 8'hca;    Blue = 8'h4a;
end 13'h7fa:    begin Red = 8'h8f;    Green = 8'h84;    Blue = 8'h61;
end 13'h7fb:    begin Red = 8'h6d;    Green = 8'h84;    Blue = 8'h42;
end 13'h7fc:    begin Red = 8'hc1;    Green = 8'had;    Blue = 8'h95;
end 13'h7fd:    begin Red = 8'hc3;    Green = 8'h8c;    Blue = 8'hb9;
end 13'h7fe:    begin Red = 8'hbd;    Green = 8'h7d;    Blue = 8'ha7;
end 13'h7ff:    begin Red = 8'hd2;    Green = 8'he0;    Blue = 8'hd1;
end 13'h800:    begin Red = 8'hd2;    Green = 8'heb;    Blue = 8'hda;
end 13'h801:    begin Red = 8'hce;    Green = 8'ha0;    Blue = 8'hd0;
end 13'h802:    begin Red = 8'hec;    Green = 8'he5;    Blue = 8'hc8;
end 13'h803:    begin Red = 8'hdf;    Green = 8'hdb;    Blue = 8'hbd;
end 13'h804:    begin Red = 8'hf7;    Green = 8'hf3;    Blue = 8'hd2;
end 13'h805:    begin Red = 8'h9b;    Green = 8'hb9;    Blue = 8'h9f;
end 13'h806:    begin Red = 8'hb0;    Green = 8'ha6;    Blue = 8'h3e;
end 13'h807:    begin Red = 8'h8b;    Green = 8'h9c;    Blue = 8'h92;
end 13'h808:    begin Red = 8'h90;    Green = 8'ha1;    Blue = 8'h87;
end 13'h809:    begin Red = 8'h73;    Green = 8'h71;    Blue = 8'h65;
end 13'h80a:    begin Red = 8'h8a;    Green = 8'h96;    Blue = 8'h54;
end 13'h80b:    begin Red = 8'haf;    Green = 8'haa;    Blue = 8'h51;
end 13'h80c:    begin Red = 8'hac;    Green = 8'ha4;    Blue = 8'h4a;
end 13'h80d:    begin Red = 8'ha7;    Green = 8'ha4;    Blue = 8'h49;
end 13'h80e:    begin Red = 8'he0;    Green = 8'hb6;    Blue = 8'h93;
end 13'h80f:    begin Red = 8'hc5;    Green = 8'hc5;    Blue = 8'h4f;
end 13'h810:    begin Red = 8'h59;    Green = 8'h6f;    Blue = 8'h41;
end 13'h811:    begin Red = 8'hb2;    Green = 8'ha1;    Blue = 8'h57;
end 13'h812:    begin Red = 8'ha1;    Green = 8'ha7;    Blue = 8'h52;
end 13'h813:    begin Red = 8'hd3;    Green = 8'hce;    Blue = 8'h5f;
end 13'h814:    begin Red = 8'hbe;    Green = 8'hd9;    Blue = 8'h54;
end 13'h815:    begin Red = 8'ha1;    Green = 8'hbb;    Blue = 8'h4d;
end 13'h816:    begin Red = 8'h69;    Green = 8'h61;    Blue = 8'h55;
end 13'h817:    begin Red = 8'ha5;    Green = 8'hc2;    Blue = 8'h44;
end 13'h818:    begin Red = 8'ha3;    Green = 8'hc0;    Blue = 8'h43;
end 13'h819:    begin Red = 8'ha2;    Green = 8'h86;    Blue = 8'h5a;
end 13'h81a:    begin Red = 8'h66;    Green = 8'h5f;    Blue = 8'h46;
end 13'h81b:    begin Red = 8'h5d;    Green = 8'h57;    Blue = 8'h45;
end 13'h81c:    begin Red = 8'h80;    Green = 8'h73;    Blue = 8'h4a;
end 13'h81d:    begin Red = 8'h7f;    Green = 8'h75;    Blue = 8'h47;
end 13'h81e:    begin Red = 8'h7d;    Green = 8'h73;    Blue = 8'h45;
end 13'h81f:    begin Red = 8'h9e;    Green = 8'h73;    Blue = 8'h4e;
end 13'h820:    begin Red = 8'h99;    Green = 8'h76;    Blue = 8'h51;
end 13'h821:    begin Red = 8'hea;    Green = 8'hd3;    Blue = 8'had;
end 13'h822:    begin Red = 8'h78;    Green = 8'h6c;    Blue = 8'h5f;
end 13'h823:    begin Red = 8'ha2;    Green = 8'h90;    Blue = 8'h66;
end 13'h824:    begin Red = 8'hd7;    Green = 8'hcb;    Blue = 8'h5a;
end 13'h825:    begin Red = 8'hcd;    Green = 8'hbd;    Blue = 8'h5a;
end 13'h826:    begin Red = 8'h9c;    Green = 8'h9b;    Blue = 8'h57;
end 13'h827:    begin Red = 8'he0;    Green = 8'hd6;    Blue = 8'h61;
end 13'h828:    begin Red = 8'ha4;    Green = 8'hc0;    Blue = 8'h47;
end 13'h829:    begin Red = 8'hbe;    Green = 8'h79;    Blue = 8'hb5;
end 13'h82a:    begin Red = 8'hd8;    Green = 8'hd2;    Blue = 8'hdc;
end 13'h82b:    begin Red = 8'hd0;    Green = 8'he5;    Blue = 8'he2;
end 13'h82c:    begin Red = 8'hd1;    Green = 8'h9d;    Blue = 8'hbe;
end 13'h82d:    begin Red = 8'hdb;    Green = 8'hd6;    Blue = 8'hbb;
end 13'h82e:    begin Red = 8'hf3;    Green = 8'hef;    Blue = 8'hce;
end 13'h82f:    begin Red = 8'hce;    Green = 8'hcf;    Blue = 8'ha7;
end 13'h830:    begin Red = 8'haf;    Green = 8'h9b;    Blue = 8'h57;
end 13'h831:    begin Red = 8'h76;    Green = 8'h77;    Blue = 8'h5e;
end 13'h832:    begin Red = 8'hc2;    Green = 8'hc1;    Blue = 8'h4e;
end 13'h833:    begin Red = 8'h63;    Green = 8'h5d;    Blue = 8'h4e;
end 13'h834:    begin Red = 8'h75;    Green = 8'h6d;    Blue = 8'h56;
end 13'h835:    begin Red = 8'hb9;    Green = 8'hd4;    Blue = 8'h42;
end 13'h836:    begin Red = 8'hb7;    Green = 8'hd8;    Blue = 8'h42;
end 13'h837:    begin Red = 8'h69;    Green = 8'h68;    Blue = 8'h57;
end 13'h838:    begin Red = 8'ha0;    Green = 8'hbe;    Blue = 8'h41;
end 13'h839:    begin Red = 8'h6f;    Green = 8'h66;    Blue = 8'h50;
end 13'h83a:    begin Red = 8'h90;    Green = 8'h82;    Blue = 8'h5f;
end 13'h83b:    begin Red = 8'h76;    Green = 8'h79;    Blue = 8'h4a;
end 13'h83c:    begin Red = 8'hab;    Green = 8'h88;    Blue = 8'h5d;
end 13'h83d:    begin Red = 8'h80;    Green = 8'h76;    Blue = 8'h50;
end 13'h83e:    begin Red = 8'h64;    Green = 8'h71;    Blue = 8'h54;
end 13'h83f:    begin Red = 8'hc8;    Green = 8'hc2;    Blue = 8'ha5;
end 13'h840:    begin Red = 8'h7e;    Green = 8'h77;    Blue = 8'h4b;
end 13'h841:    begin Red = 8'h7c;    Green = 8'h75;    Blue = 8'h49;
end 13'h842:    begin Red = 8'hfd;    Green = 8'heb;    Blue = 8'hc6;
end 13'h843:    begin Red = 8'hef;    Green = 8'hdd;    Blue = 8'hbb;
end 13'h844:    begin Red = 8'h88;    Green = 8'h7b;    Blue = 8'h6b;
end 13'h845:    begin Red = 8'h9a;    Green = 8'h8b;    Blue = 8'h73;
end 13'h846:    begin Red = 8'hfd;    Green = 8'he4;    Blue = 8'hd3;
end 13'h847:    begin Red = 8'hff;    Green = 8'hf1;    Blue = 8'he6;
end 13'h848:    begin Red = 8'hcc;    Green = 8'hc7;    Blue = 8'h5b;
end 13'h849:    begin Red = 8'h5b;    Green = 8'h69;    Blue = 8'h4c;
end 13'h84a:    begin Red = 8'h51;    Green = 8'h49;    Blue = 8'h42;
end 13'h84b:    begin Red = 8'h59;    Green = 8'h4e;    Blue = 8'h45;
end 13'h84c:    begin Red = 8'h8e;    Green = 8'h83;    Blue = 8'h5c;
end 13'h84d:    begin Red = 8'h5f;    Green = 8'h58;    Blue = 8'h52;
end 13'h84e:    begin Red = 8'h92;    Green = 8'h80;    Blue = 8'h5e;
end 13'h84f:    begin Red = 8'h5e;    Green = 8'h5a;    Blue = 8'h57;
end 13'h850:    begin Red = 8'h93;    Green = 8'ha0;    Blue = 8'h62;
end 13'h851:    begin Red = 8'hc3;    Green = 8'hcc;    Blue = 8'hc7;
end 13'h852:    begin Red = 8'hb2;    Green = 8'hcc;    Blue = 8'hb5;
end 13'h853:    begin Red = 8'hd6;    Green = 8'h91;    Blue = 8'hc8;
end 13'h854:    begin Red = 8'hce;    Green = 8'h8e;    Blue = 8'hbd;
end 13'h855:    begin Red = 8'hd8;    Green = 8'hd5;    Blue = 8'hb9;
end 13'h856:    begin Red = 8'hf2;    Green = 8'he8;    Blue = 8'hbe;
end 13'h857:    begin Red = 8'hac;    Green = 8'ha5;    Blue = 8'h45;
end 13'h858:    begin Red = 8'hb0;    Green = 8'ha4;    Blue = 8'h52;
end 13'h859:    begin Red = 8'hb5;    Green = 8'hcb;    Blue = 8'h42;
end 13'h85a:    begin Red = 8'h61;    Green = 8'h61;    Blue = 8'h58;
end 13'h85b:    begin Red = 8'ha7;    Green = 8'hbb;    Blue = 8'h43;
end 13'h85c:    begin Red = 8'h85;    Green = 8'h8b;    Blue = 8'h61;
end 13'h85d:    begin Red = 8'hde;    Green = 8'hb1;    Blue = 8'h94;
end 13'h85e:    begin Red = 8'h8e;    Green = 8'h6c;    Blue = 8'h65;
end 13'h85f:    begin Red = 8'ha0;    Green = 8'h7b;    Blue = 8'h71;
end 13'h860:    begin Red = 8'hd3;    Green = 8'hca;    Blue = 8'h53;
end 13'h861:    begin Red = 8'h51;    Green = 8'h66;    Blue = 8'h42;
end 13'h862:    begin Red = 8'h53;    Green = 8'h48;    Blue = 8'h3f;
end 13'h863:    begin Red = 8'h6b;    Green = 8'h61;    Blue = 8'h3f;
end 13'h864:    begin Red = 8'h90;    Green = 8'h82;    Blue = 8'h5a;
end 13'h865:    begin Red = 8'h65;    Green = 8'h55;    Blue = 8'h59;
end 13'h866:    begin Red = 8'h67;    Green = 8'h5a;    Blue = 8'h50;
end 13'h867:    begin Red = 8'h89;    Green = 8'h96;    Blue = 8'h5d;
end 13'h868:    begin Red = 8'h9e;    Green = 8'h82;    Blue = 8'h4f;
end 13'h869:    begin Red = 8'haf;    Green = 8'h88;    Blue = 8'h57;
end 13'h86a:    begin Red = 8'h62;    Green = 8'h66;    Blue = 8'h4e;
end 13'h86b:    begin Red = 8'haf;    Green = 8'haf;    Blue = 8'h93;
end 13'h86c:    begin Red = 8'h82;    Green = 8'h74;    Blue = 8'h57;
end 13'h86d:    begin Red = 8'h87;    Green = 8'h75;    Blue = 8'h4b;
end 13'h86e:    begin Red = 8'h81;    Green = 8'h73;    Blue = 8'h60;
end 13'h86f:    begin Red = 8'hf3;    Green = 8'he2;    Blue = 8'hb7;
end 13'h870:    begin Red = 8'hbd;    Green = 8'hbb;    Blue = 8'h52;
end 13'h871:    begin Red = 8'hb6;    Green = 8'haa;    Blue = 8'h5a;
end 13'h872:    begin Red = 8'h62;    Green = 8'h5a;    Blue = 8'h3e;
end 13'h873:    begin Red = 8'h86;    Green = 8'h7e;    Blue = 8'h55;
end 13'h874:    begin Red = 8'h84;    Green = 8'h7d;    Blue = 8'h5b;
end 13'h875:    begin Red = 8'h65;    Green = 8'h63;    Blue = 8'h3f;
end 13'h876:    begin Red = 8'h6c;    Green = 8'h78;    Blue = 8'h4f;
end 13'h877:    begin Red = 8'hb8;    Green = 8'hc2;    Blue = 8'hb2;
end 13'h878:    begin Red = 8'hd9;    Green = 8'h9e;    Blue = 8'hca;
end 13'h879:    begin Red = 8'hd6;    Green = 8'h9c;    Blue = 8'hc3;
end 13'h87a:    begin Red = 8'hd8;    Green = 8'h98;    Blue = 8'hc7;
end 13'h87b:    begin Red = 8'hf6;    Green = 8'hf1;    Blue = 8'hcf;
end 13'h87c:    begin Red = 8'hfd;    Green = 8'hf7;    Blue = 8'hd6;
end 13'h87d:    begin Red = 8'ha3;    Green = 8'haf;    Blue = 8'h9f;
end 13'h87e:    begin Red = 8'h8a;    Green = 8'h86;    Blue = 8'h68;
end 13'h87f:    begin Red = 8'h94;    Green = 8'h7a;    Blue = 8'h5a;
end 13'h880:    begin Red = 8'h61;    Green = 8'h61;    Blue = 8'h4d;
end 13'h881:    begin Red = 8'ha4;    Green = 8'h84;    Blue = 8'h59;
end 13'h882:    begin Red = 8'h88;    Green = 8'h76;    Blue = 8'h55;
end 13'h883:    begin Red = 8'h6e;    Green = 8'h77;    Blue = 8'h5c;
end 13'h884:    begin Red = 8'hb6;    Green = 8'haf;    Blue = 8'h94;
end 13'h885:    begin Red = 8'ha2;    Green = 8'h9f;    Blue = 8'h80;
end 13'h886:    begin Red = 8'haa;    Green = 8'hab;    Blue = 8'h92;
end 13'h887:    begin Red = 8'h9a;    Green = 8'h7d;    Blue = 8'h4f;
end 13'h888:    begin Red = 8'hd7;    Green = 8'hc7;    Blue = 8'ha3;
end 13'h889:    begin Red = 8'h52;    Green = 8'h55;    Blue = 8'h3b;
end 13'h88a:    begin Red = 8'h67;    Green = 8'h5d;    Blue = 8'h49;
end 13'h88b:    begin Red = 8'hb8;    Green = 8'h98;    Blue = 8'h69;
end 13'h88c:    begin Red = 8'hcf;    Green = 8'hd7;    Blue = 8'hd8;
end 13'h88d:    begin Red = 8'hd9;    Green = 8'hd7;    Blue = 8'he0;
end 13'h88e:    begin Red = 8'hd7;    Green = 8'hd2;    Blue = 8'hb0;
end 13'h88f:    begin Red = 8'h7d;    Green = 8'h86;    Blue = 8'h60;
end 13'h890:    begin Red = 8'ha3;    Green = 8'hbb;    Blue = 8'h42;
end 13'h891:    begin Red = 8'h88;    Green = 8'h98;    Blue = 8'h94;
end 13'h892:    begin Red = 8'h6f;    Green = 8'h8d;    Blue = 8'h4a;
end 13'h893:    begin Red = 8'h6c;    Green = 8'h62;    Blue = 8'h44;
end 13'h894:    begin Red = 8'hb7;    Green = 8'h92;    Blue = 8'h6a;
end 13'h895:    begin Red = 8'hb8;    Green = 8'h90;    Blue = 8'h6d;
end 13'h896:    begin Red = 8'h5d;    Green = 8'h59;    Blue = 8'h3c;
end 13'h897:    begin Red = 8'h69;    Green = 8'h62;    Blue = 8'h4a;
end 13'h898:    begin Red = 8'hf1;    Green = 8'hf1;    Blue = 8'hc6;
end 13'h899:    begin Red = 8'hcf;    Green = 8'hca;    Blue = 8'hb3;
end 13'h89a:    begin Red = 8'hb1;    Green = 8'h89;    Blue = 8'h5a;
end 13'h89b:    begin Red = 8'h66;    Green = 8'h6e;    Blue = 8'h5a;
end 13'h89c:    begin Red = 8'h60;    Green = 8'h67;    Blue = 8'h51;
end 13'h89d:    begin Red = 8'ha3;    Green = 8'h9f;    Blue = 8'h85;
end 13'h89e:    begin Red = 8'ha5;    Green = 8'ha4;    Blue = 8'h8c;
end 13'h89f:    begin Red = 8'hfd;    Green = 8'heb;    Blue = 8'hcc;
end 13'h8a0:    begin Red = 8'ha3;    Green = 8'h7b;    Blue = 8'h4f;
end 13'h8a1:    begin Red = 8'h7d;    Green = 8'h6f;    Blue = 8'h5d;
end 13'h8a2:    begin Red = 8'h7f;    Green = 8'h74;    Blue = 8'h5e;
end 13'h8a3:    begin Red = 8'h62;    Green = 8'h7e;    Blue = 8'h3d;
end 13'h8a4:    begin Red = 8'h76;    Green = 8'h93;    Blue = 8'h4b;
end 13'h8a5:    begin Red = 8'h86;    Green = 8'h75;    Blue = 8'h4f;
end 13'h8a6:    begin Red = 8'h65;    Green = 8'h61;    Blue = 8'h3a;
end 13'h8a7:    begin Red = 8'hcf;    Green = 8'ha0;    Blue = 8'h76;
end 13'h8a8:    begin Red = 8'hbf;    Green = 8'ha0;    Blue = 8'h71;
end 13'h8a9:    begin Red = 8'hc3;    Green = 8'h9e;    Blue = 8'h75;
end 13'h8aa:    begin Red = 8'hbe;    Green = 8'h93;    Blue = 8'h6e;
end 13'h8ab:    begin Red = 8'h85;    Green = 8'h9c;    Blue = 8'h5b;
end 13'h8ac:    begin Red = 8'h7a;    Green = 8'h94;    Blue = 8'h57;
end 13'h8ad:    begin Red = 8'hba;    Green = 8'hc3;    Blue = 8'hc6;
end 13'h8ae:    begin Red = 8'hd5;    Green = 8'h96;    Blue = 8'hc3;
end 13'h8af:    begin Red = 8'hd7;    Green = 8'h95;    Blue = 8'hce;
end 13'h8b0:    begin Red = 8'hd3;    Green = 8'h8c;    Blue = 8'hce;
end 13'h8b1:    begin Red = 8'hff;    Green = 8'hfa;    Blue = 8'hd7;
end 13'h8b2:    begin Red = 8'he4;    Green = 8'hda;    Blue = 8'hb9;
end 13'h8b3:    begin Red = 8'hf3;    Green = 8'he5;    Blue = 8'hc0;
end 13'h8b4:    begin Red = 8'h79;    Green = 8'h89;    Blue = 8'h75;
end 13'h8b5:    begin Red = 8'h9b;    Green = 8'hb6;    Blue = 8'h8e;
end 13'h8b6:    begin Red = 8'h94;    Green = 8'hb9;    Blue = 8'ha9;
end 13'h8b7:    begin Red = 8'hc8;    Green = 8'hc5;    Blue = 8'h61;
end 13'h8b8:    begin Red = 8'hb7;    Green = 8'hd7;    Blue = 8'h46;
end 13'h8b9:    begin Red = 8'hb0;    Green = 8'hce;    Blue = 8'h45;
end 13'h8ba:    begin Red = 8'ha2;    Green = 8'hb5;    Blue = 8'h46;
end 13'h8bb:    begin Red = 8'h79;    Green = 8'h98;    Blue = 8'h85;
end 13'h8bc:    begin Red = 8'h65;    Green = 8'h82;    Blue = 8'h42;
end 13'h8bd:    begin Red = 8'h7f;    Green = 8'h90;    Blue = 8'h54;
end 13'h8be:    begin Red = 8'h79;    Green = 8'h87;    Blue = 8'h5b;
end 13'h8bf:    begin Red = 8'h8c;    Green = 8'h7d;    Blue = 8'h50;
end 13'h8c0:    begin Red = 8'h53;    Green = 8'h53;    Blue = 8'h3d;
end 13'h8c1:    begin Red = 8'hbf;    Green = 8'ha2;    Blue = 8'h78;
end 13'h8c2:    begin Red = 8'h8f;    Green = 8'h7d;    Blue = 8'h5a;
end 13'h8c3:    begin Red = 8'hbc;    Green = 8'h96;    Blue = 8'h71;
end 13'h8c4:    begin Red = 8'h7b;    Green = 8'h7d;    Blue = 8'h55;
end 13'h8c5:    begin Red = 8'hf7;    Green = 8'hc3;    Blue = 8'h95;
end 13'h8c6:    begin Red = 8'hfb;    Green = 8'hcc;    Blue = 8'ha0;
end 13'h8c7:    begin Red = 8'he4;    Green = 8'hdc;    Blue = 8'hb2;
end 13'h8c8:    begin Red = 8'he9;    Green = 8'he2;    Blue = 8'hb6;
end 13'h8c9:    begin Red = 8'hc3;    Green = 8'hbc;    Blue = 8'h9b;
end 13'h8ca:    begin Red = 8'h9d;    Green = 8'h83;    Blue = 8'h59;
end 13'h8cb:    begin Red = 8'h6c;    Green = 8'h76;    Blue = 8'h56;
end 13'h8cc:    begin Red = 8'ha2;    Green = 8'ha9;    Blue = 8'h98;
end 13'h8cd:    begin Red = 8'ha0;    Green = 8'h7d;    Blue = 8'h4f;
end 13'h8ce:    begin Red = 8'h82;    Green = 8'h79;    Blue = 8'h46;
end 13'h8cf:    begin Red = 8'h72;    Green = 8'h85;    Blue = 8'h42;
end 13'h8d0:    begin Red = 8'hc3;    Green = 8'ha2;    Blue = 8'h72;
end 13'h8d1:    begin Red = 8'had;    Green = 8'h92;    Blue = 8'h6d;
end 13'h8d2:    begin Red = 8'h7d;    Green = 8'h7c;    Blue = 8'h51;
end 13'h8d3:    begin Red = 8'hb7;    Green = 8'h99;    Blue = 8'h6f;
end 13'h8d4:    begin Red = 8'h69;    Green = 8'h61;    Blue = 8'h45;
end 13'h8d5:    begin Red = 8'hd0;    Green = 8'hbe;    Blue = 8'h9c;
end 13'h8d6:    begin Red = 8'hba;    Green = 8'hc0;    Blue = 8'hc3;
end 13'h8d7:    begin Red = 8'hbe;    Green = 8'hbb;    Blue = 8'hc0;
end 13'h8d8:    begin Red = 8'hd2;    Green = 8'ha0;    Blue = 8'hd8;
end 13'h8d9:    begin Red = 8'hd9;    Green = 8'h9b;    Blue = 8'hc1;
end 13'h8da:    begin Red = 8'hda;    Green = 8'h8f;    Blue = 8'hbd;
end 13'h8db:    begin Red = 8'hd4;    Green = 8'hd0;    Blue = 8'haf;
end 13'h8dc:    begin Red = 8'hb3;    Green = 8'ha8;    Blue = 8'h57;
end 13'h8dd:    begin Red = 8'ha8;    Green = 8'hbf;    Blue = 8'h50;
end 13'h8de:    begin Red = 8'h80;    Green = 8'h90;    Blue = 8'h59;
end 13'h8df:    begin Red = 8'h80;    Green = 8'h8f;    Blue = 8'h9a;
end 13'h8e0:    begin Red = 8'hdf;    Green = 8'hb1;    Blue = 8'h8c;
end 13'h8e1:    begin Red = 8'h54;    Green = 8'h50;    Blue = 8'h39;
end 13'h8e2:    begin Red = 8'hb3;    Green = 8'h92;    Blue = 8'h6c;
end 13'h8e3:    begin Red = 8'h7a;    Green = 8'h7a;    Blue = 8'h52;
end 13'h8e4:    begin Red = 8'h8c;    Green = 8'h7c;    Blue = 8'h56;
end 13'h8e5:    begin Red = 8'h8c;    Green = 8'h79;    Blue = 8'h5e;
end 13'h8e6:    begin Red = 8'h7c;    Green = 8'h7b;    Blue = 8'h58;
end 13'h8e7:    begin Red = 8'hb5;    Green = 8'h93;    Blue = 8'h67;
end 13'h8e8:    begin Red = 8'hc6;    Green = 8'hbb;    Blue = 8'ha0;
end 13'h8e9:    begin Red = 8'h9c;    Green = 8'ha5;    Blue = 8'h75;
end 13'h8ea:    begin Red = 8'h92;    Green = 8'h9b;    Blue = 8'h78;
end 13'h8eb:    begin Red = 8'h8e;    Green = 8'h94;    Blue = 8'h6d;
end 13'h8ec:    begin Red = 8'h97;    Green = 8'h70;    Blue = 8'h42;
end 13'h8ed:    begin Red = 8'h99;    Green = 8'h71;    Blue = 8'h4b;
end 13'h8ee:    begin Red = 8'ha5;    Green = 8'h8d;    Blue = 8'h6f;
end 13'h8ef:    begin Red = 8'h88;    Green = 8'h7c;    Blue = 8'h46;
end 13'h8f0:    begin Red = 8'h86;    Green = 8'h7d;    Blue = 8'h51;
end 13'h8f1:    begin Red = 8'h62;    Green = 8'h60;    Blue = 8'h3f;
end 13'h8f2:    begin Red = 8'haf;    Green = 8'h92;    Blue = 8'h71;
end 13'h8f3:    begin Red = 8'h69;    Green = 8'h5c;    Blue = 8'h47;
end 13'h8f4:    begin Red = 8'h7f;    Green = 8'h76;    Blue = 8'h42;
end 13'h8f5:    begin Red = 8'hc5;    Green = 8'hbb;    Blue = 8'hca;
end 13'h8f6:    begin Red = 8'hc9;    Green = 8'h91;    Blue = 8'hbb;
end 13'h8f7:    begin Red = 8'hc4;    Green = 8'h83;    Blue = 8'hb4;
end 13'h8f8:    begin Red = 8'hdb;    Green = 8'ha0;    Blue = 8'hc9;
end 13'h8f9:    begin Red = 8'ha0;    Green = 8'hb5;    Blue = 8'h8c;
end 13'h8fa:    begin Red = 8'h8b;    Green = 8'hb5;    Blue = 8'ha8;
end 13'h8fb:    begin Red = 8'h9d;    Green = 8'ha3;    Blue = 8'h51;
end 13'h8fc:    begin Red = 8'h95;    Green = 8'ha8;    Blue = 8'h4f;
end 13'h8fd:    begin Red = 8'h8c;    Green = 8'h89;    Blue = 8'h5d;
end 13'h8fe:    begin Red = 8'h5b;    Green = 8'h58;    Blue = 8'h41;
end 13'h8ff:    begin Red = 8'h84;    Green = 8'h77;    Blue = 8'h48;
end 13'h900:    begin Red = 8'h71;    Green = 8'h63;    Blue = 8'h3f;
end 13'h901:    begin Red = 8'hd6;    Green = 8'hb3;    Blue = 8'h82;
end 13'h902:    begin Red = 8'hd5;    Green = 8'hb0;    Blue = 8'h87;
end 13'h903:    begin Red = 8'hc4;    Green = 8'hbe;    Blue = 8'ha0;
end 13'h904:    begin Red = 8'h9d;    Green = 8'ha0;    Blue = 8'h78;
end 13'h905:    begin Red = 8'h9e;    Green = 8'ha5;    Blue = 8'h78;
end 13'h906:    begin Red = 8'h90;    Green = 8'h95;    Blue = 8'h77;
end 13'h907:    begin Red = 8'h64;    Green = 8'h69;    Blue = 8'h52;
end 13'h908:    begin Red = 8'h8b;    Green = 8'h5e;    Blue = 8'h34;
end 13'h909:    begin Red = 8'h84;    Green = 8'h64;    Blue = 8'h3f;
end 13'h90a:    begin Red = 8'h8e;    Green = 8'h66;    Blue = 8'h37;
end 13'h90b:    begin Red = 8'h8c;    Green = 8'h66;    Blue = 8'h42;
end 13'h90c:    begin Red = 8'hec;    Green = 8'hd6;    Blue = 8'hb6;
end 13'h90d:    begin Red = 8'haf;    Green = 8'h9b;    Blue = 8'h87;
end 13'h90e:    begin Red = 8'hb0;    Green = 8'h96;    Blue = 8'h8a;
end 13'h90f:    begin Red = 8'h7d;    Green = 8'h71;    Blue = 8'h4c;
end 13'h910:    begin Red = 8'h7d;    Green = 8'h81;    Blue = 8'h56;
end 13'h911:    begin Red = 8'hc2;    Green = 8'h9a;    Blue = 8'h70;
end 13'h912:    begin Red = 8'h84;    Green = 8'h72;    Blue = 8'h44;
end 13'h913:    begin Red = 8'h81;    Green = 8'h72;    Blue = 8'h46;
end 13'h914:    begin Red = 8'hb0;    Green = 8'h97;    Blue = 8'h83;
end 13'h915:    begin Red = 8'hf9;    Green = 8'hce;    Blue = 8'hb3;
end 13'h916:    begin Red = 8'h79;    Green = 8'h96;    Blue = 8'h4e;
end 13'h917:    begin Red = 8'h70;    Green = 8'h83;    Blue = 8'h3d;
end 13'h918:    begin Red = 8'h71;    Green = 8'h88;    Blue = 8'h47;
end 13'h919:    begin Red = 8'h66;    Green = 8'h90;    Blue = 8'h4a;
end 13'h91a:    begin Red = 8'h8a;    Green = 8'h77;    Blue = 8'h61;
end 13'h91b:    begin Red = 8'hc2;    Green = 8'h84;    Blue = 8'hac;
end 13'h91c:    begin Red = 8'hd7;    Green = 8'hd9;    Blue = 8'hcc;
end 13'h91d:    begin Red = 8'hd1;    Green = 8'hec;    Blue = 8'hdf;
end 13'h91e:    begin Red = 8'hd8;    Green = 8'ha3;    Blue = 8'hcb;
end 13'h91f:    begin Red = 8'hd2;    Green = 8'hdf;    Blue = 8'hd7;
end 13'h920:    begin Red = 8'hc6;    Green = 8'hc0;    Blue = 8'h9f;
end 13'h921:    begin Red = 8'hd0;    Green = 8'hca;    Blue = 8'ha9;
end 13'h922:    begin Red = 8'h71;    Green = 8'h88;    Blue = 8'h78;
end 13'h923:    begin Red = 8'h98;    Green = 8'hb3;    Blue = 8'ha6;
end 13'h924:    begin Red = 8'h9a;    Green = 8'h96;    Blue = 8'h46;
end 13'h925:    begin Red = 8'h82;    Green = 8'h87;    Blue = 8'h64;
end 13'h926:    begin Red = 8'h80;    Green = 8'h8f;    Blue = 8'h4c;
end 13'h927:    begin Red = 8'h9f;    Green = 8'hb7;    Blue = 8'h37;
end 13'h928:    begin Red = 8'h78;    Green = 8'h80;    Blue = 8'h65;
end 13'h929:    begin Red = 8'h94;    Green = 8'ha8;    Blue = 8'h41;
end 13'h92a:    begin Red = 8'h84;    Green = 8'h9d;    Blue = 8'h8c;
end 13'h92b:    begin Red = 8'h78;    Green = 8'h9b;    Blue = 8'h89;
end 13'h92c:    begin Red = 8'hac;    Green = 8'h98;    Blue = 8'h77;
end 13'h92d:    begin Red = 8'h5d;    Green = 8'h5a;    Blue = 8'h42;
end 13'h92e:    begin Red = 8'h94;    Green = 8'h8f;    Blue = 8'h64;
end 13'h92f:    begin Red = 8'h8a;    Green = 8'h88;    Blue = 8'h65;
end 13'h930:    begin Red = 8'h7f;    Green = 8'h77;    Blue = 8'h5b;
end 13'h931:    begin Red = 8'hc2;    Green = 8'h90;    Blue = 8'h73;
end 13'h932:    begin Red = 8'h55;    Green = 8'h55;    Blue = 8'h39;
end 13'h933:    begin Red = 8'h8b;    Green = 8'h82;    Blue = 8'h5e;
end 13'h934:    begin Red = 8'h65;    Green = 8'h5f;    Blue = 8'h3e;
end 13'h935:    begin Red = 8'h75;    Green = 8'h71;    Blue = 8'h3c;
end 13'h936:    begin Red = 8'hed;    Green = 8'hc3;    Blue = 8'h9a;
end 13'h937:    begin Red = 8'h9a;    Green = 8'ha1;    Blue = 8'h75;
end 13'h938:    begin Red = 8'heb;    Green = 8'hd9;    Blue = 8'hb8;
end 13'h939:    begin Red = 8'h90;    Green = 8'h7d;    Blue = 8'h66;
end 13'h93a:    begin Red = 8'h8f;    Green = 8'h7a;    Blue = 8'h65;
end 13'h93b:    begin Red = 8'hb2;    Green = 8'h98;    Blue = 8'h8e;
end 13'h93c:    begin Red = 8'haa;    Green = 8'h87;    Blue = 8'h55;
end 13'h93d:    begin Red = 8'h63;    Green = 8'h55;    Blue = 8'h42;
end 13'h93e:    begin Red = 8'hc5;    Green = 8'h9c;    Blue = 8'h72;
end 13'h93f:    begin Red = 8'h89;    Green = 8'h78;    Blue = 8'h4d;
end 13'h940:    begin Red = 8'h90;    Green = 8'h74;    Blue = 8'h61;
end 13'h941:    begin Red = 8'h8e;    Green = 8'h7a;    Blue = 8'h61;
end 13'h942:    begin Red = 8'hca;    Green = 8'h93;    Blue = 8'hbe;
end 13'h943:    begin Red = 8'hd6;    Green = 8'ha3;    Blue = 8'hc7;
end 13'h944:    begin Red = 8'hda;    Green = 8'ha6;    Blue = 8'hcc;
end 13'h945:    begin Red = 8'hd2;    Green = 8'h9f;    Blue = 8'hcd;
end 13'h946:    begin Red = 8'heb;    Green = 8'he9;    Blue = 8'hc8;
end 13'h947:    begin Red = 8'hf9;    Green = 8'hf6;    Blue = 8'hd2;
end 13'h948:    begin Red = 8'h72;    Green = 8'h86;    Blue = 8'h75;
end 13'h949:    begin Red = 8'h98;    Green = 8'hb4;    Blue = 8'h9b;
end 13'h94a:    begin Red = 8'h9e;    Green = 8'hbb;    Blue = 8'haf;
end 13'h94b:    begin Red = 8'ha6;    Green = 8'ha7;    Blue = 8'h52;
end 13'h94c:    begin Red = 8'h7d;    Green = 8'h78;    Blue = 8'h6b;
end 13'h94d:    begin Red = 8'h46;    Green = 8'h4b;    Blue = 8'h42;
end 13'h94e:    begin Red = 8'h74;    Green = 8'h7a;    Blue = 8'h55;
end 13'h94f:    begin Red = 8'h97;    Green = 8'ha9;    Blue = 8'h53;
end 13'h950:    begin Red = 8'ha9;    Green = 8'h82;    Blue = 8'h55;
end 13'h951:    begin Red = 8'hb4;    Green = 8'h8f;    Blue = 8'h6d;
end 13'h952:    begin Red = 8'h8a;    Green = 8'h7b;    Blue = 8'h4c;
end 13'h953:    begin Red = 8'hed;    Green = 8'hc3;    Blue = 8'ha0;
end 13'h954:    begin Red = 8'h8f;    Green = 8'h94;    Blue = 8'h74;
end 13'h955:    begin Red = 8'hb7;    Green = 8'h99;    Blue = 8'h7d;
end 13'h956:    begin Red = 8'h9c;    Green = 8'h84;    Blue = 8'h6d;
end 13'h957:    begin Red = 8'h82;    Green = 8'h9b;    Blue = 8'h3a;
end 13'h958:    begin Red = 8'hf1;    Green = 8'hdf;    Blue = 8'hb6;
end 13'h959:    begin Red = 8'h81;    Green = 8'h9e;    Blue = 8'h35;
end 13'h95a:    begin Red = 8'h98;    Green = 8'ha4;    Blue = 8'h43;
end 13'h95b:    begin Red = 8'h92;    Green = 8'ha7;    Blue = 8'h52;
end 13'h95c:    begin Red = 8'h7e;    Green = 8'h78;    Blue = 8'h51;
end 13'h95d:    begin Red = 8'ha6;    Green = 8'h86;    Blue = 8'h57;
end 13'h95e:    begin Red = 8'h56;    Green = 8'h58;    Blue = 8'h46;
end 13'h95f:    begin Red = 8'h87;    Green = 8'h7d;    Blue = 8'h4d;
end 13'h960:    begin Red = 8'hd0;    Green = 8'he2;    Blue = 8'hd7;
end 13'h961:    begin Red = 8'hd6;    Green = 8'ha3;    Blue = 8'hce;
end 13'h962:    begin Red = 8'hb9;    Green = 8'hb6;    Blue = 8'h9f;
end 13'h963:    begin Red = 8'hc1;    Green = 8'hbd;    Blue = 8'ha5;
end 13'h964:    begin Red = 8'hc4;    Green = 8'hc1;    Blue = 8'ha5;
end 13'h965:    begin Red = 8'hd3;    Green = 8'hce;    Blue = 8'hb2;
end 13'h966:    begin Red = 8'hb5;    Green = 8'hb2;    Blue = 8'h96;
end 13'h967:    begin Red = 8'hb6;    Green = 8'hb2;    Blue = 8'ha0;
end 13'h968:    begin Red = 8'hb4;    Green = 8'hb1;    Blue = 8'h9b;
end 13'h969:    begin Red = 8'hce;    Green = 8'hc4;    Blue = 8'h4e;
end 13'h96a:    begin Red = 8'hb5;    Green = 8'hce;    Blue = 8'h4a;
end 13'h96b:    begin Red = 8'hac;    Green = 8'hc6;    Blue = 8'h4f;
end 13'h96c:    begin Red = 8'hba;    Green = 8'hcf;    Blue = 8'h44;
end 13'h96d:    begin Red = 8'h43;    Green = 8'h4d;    Blue = 8'h43;
end 13'h96e:    begin Red = 8'h87;    Green = 8'ha3;    Blue = 8'h43;
end 13'h96f:    begin Red = 8'h84;    Green = 8'ha8;    Blue = 8'h4a;
end 13'h970:    begin Red = 8'ha6;    Green = 8'h7c;    Blue = 8'h63;
end 13'h971:    begin Red = 8'ha3;    Green = 8'h7b;    Blue = 8'h6a;
end 13'h972:    begin Red = 8'h94;    Green = 8'had;    Blue = 8'h48;
end 13'h973:    begin Red = 8'h84;    Green = 8'haf;    Blue = 8'h92;
end 13'h974:    begin Red = 8'h94;    Green = 8'haa;    Blue = 8'h52;
end 13'h975:    begin Red = 8'h88;    Green = 8'h72;    Blue = 8'h48;
end 13'h976:    begin Red = 8'h5c;    Green = 8'h53;    Blue = 8'h43;
end 13'h977:    begin Red = 8'h5f;    Green = 8'h5b;    Blue = 8'h4a;
end 13'h978:    begin Red = 8'h94;    Green = 8'h78;    Blue = 8'h4d;
end 13'h979:    begin Red = 8'h98;    Green = 8'h75;    Blue = 8'h4e;
end 13'h97a:    begin Red = 8'h93;    Green = 8'h73;    Blue = 8'h4a;
end 13'h97b:    begin Red = 8'he5;    Green = 8'hc0;    Blue = 8'h98;
end 13'h97c:    begin Red = 8'hc2;    Green = 8'hbb;    Blue = 8'h9f;
end 13'h97d:    begin Red = 8'hab;    Green = 8'h9f;    Blue = 8'h80;
end 13'h97e:    begin Red = 8'h91;    Green = 8'had;    Blue = 8'h5d;
end 13'h97f:    begin Red = 8'hf3;    Green = 8'hdb;    Blue = 8'hbe;
end 13'h980:    begin Red = 8'h7d;    Green = 8'ha3;    Blue = 8'h3b;
end 13'h981:    begin Red = 8'hff;    Green = 8'he8;    Blue = 8'hcf;
end 13'h982:    begin Red = 8'h85;    Green = 8'h71;    Blue = 8'h53;
end 13'h983:    begin Red = 8'h98;    Green = 8'h7b;    Blue = 8'h55;
end 13'h984:    begin Red = 8'h91;    Green = 8'h7a;    Blue = 8'h4e;
end 13'h985:    begin Red = 8'he8;    Green = 8'hdd;    Blue = 8'hbf;
end 13'h986:    begin Red = 8'hc7;    Green = 8'h83;    Blue = 8'hb7;
end 13'h987:    begin Red = 8'hd0;    Green = 8'hde;    Blue = 8'hd5;
end 13'h988:    begin Red = 8'hbe;    Green = 8'hbb;    Blue = 8'ha3;
end 13'h989:    begin Red = 8'hbc;    Green = 8'hb8;    Blue = 8'h9f;
end 13'h98a:    begin Red = 8'hc6;    Green = 8'hc2;    Blue = 8'ha8;
end 13'h98b:    begin Red = 8'hb9;    Green = 8'had;    Blue = 8'h96;
end 13'h98c:    begin Red = 8'hac;    Green = 8'hb1;    Blue = 8'h93;
end 13'h98d:    begin Red = 8'h9e;    Green = 8'haf;    Blue = 8'h9f;
end 13'h98e:    begin Red = 8'hcb;    Green = 8'hc3;    Blue = 8'h50;
end 13'h98f:    begin Red = 8'h97;    Green = 8'h9a;    Blue = 8'h4d;
end 13'h990:    begin Red = 8'h83;    Green = 8'h82;    Blue = 8'h5f;
end 13'h991:    begin Red = 8'haf;    Green = 8'hc3;    Blue = 8'h4e;
end 13'h992:    begin Red = 8'hba;    Green = 8'hcd;    Blue = 8'h55;
end 13'h993:    begin Red = 8'h48;    Green = 8'h50;    Blue = 8'h3d;
end 13'h994:    begin Red = 8'h71;    Green = 8'h7a;    Blue = 8'h58;
end 13'h995:    begin Red = 8'h88;    Green = 8'ha8;    Blue = 8'h42;
end 13'h996:    begin Red = 8'hde;    Green = 8'hb8;    Blue = 8'h8d;
end 13'h997:    begin Red = 8'h8e;    Green = 8'ha5;    Blue = 8'h46;
end 13'h998:    begin Red = 8'ha0;    Green = 8'h7e;    Blue = 8'h60;
end 13'h999:    begin Red = 8'h8f;    Green = 8'hb1;    Blue = 8'h78;
end 13'h99a:    begin Red = 8'h8d;    Green = 8'haf;    Blue = 8'h83;
end 13'h99b:    begin Red = 8'h88;    Green = 8'h77;    Blue = 8'h51;
end 13'h99c:    begin Red = 8'h78;    Green = 8'h72;    Blue = 8'h4e;
end 13'h99d:    begin Red = 8'ha5;    Green = 8'h88;    Blue = 8'h59;
end 13'h99e:    begin Red = 8'h8e;    Green = 8'h7d;    Blue = 8'h4a;
end 13'h99f:    begin Red = 8'h96;    Green = 8'h73;    Blue = 8'h4c;
end 13'h9a0:    begin Red = 8'h9e;    Green = 8'ha4;    Blue = 8'h7c;
end 13'h9a1:    begin Red = 8'h7a;    Green = 8'h7e;    Blue = 8'h66;
end 13'h9a2:    begin Red = 8'h7f;    Green = 8'h84;    Blue = 8'h69;
end 13'h9a3:    begin Red = 8'h9e;    Green = 8'h94;    Blue = 8'h6e;
end 13'h9a4:    begin Red = 8'h98;    Green = 8'ha6;    Blue = 8'h4d;
end 13'h9a5:    begin Red = 8'h8d;    Green = 8'haa;    Blue = 8'h46;
end 13'h9a6:    begin Red = 8'haf;    Green = 8'ha0;    Blue = 8'h7e;
end 13'h9a7:    begin Red = 8'h9b;    Green = 8'h8f;    Blue = 8'h75;
end 13'h9a8:    begin Red = 8'h9b;    Green = 8'h8d;    Blue = 8'h80;
end 13'h9a9:    begin Red = 8'ha9;    Green = 8'h84;    Blue = 8'h5d;
end 13'h9aa:    begin Red = 8'hb2;    Green = 8'h8b;    Blue = 8'h5e;
end 13'h9ab:    begin Red = 8'h9e;    Green = 8'h87;    Blue = 8'h59;
end 13'h9ac:    begin Red = 8'h6a;    Green = 8'h77;    Blue = 8'h60;
end 13'h9ad:    begin Red = 8'h6b;    Green = 8'h5c;    Blue = 8'h34;
end 13'h9ae:    begin Red = 8'h80;    Green = 8'h7a;    Blue = 8'h48;
end 13'h9af:    begin Red = 8'h82;    Green = 8'h75;    Blue = 8'h44;
end 13'h9b0:    begin Red = 8'hf2;    Green = 8'hd9;    Blue = 8'hb0;
end 13'h9b1:    begin Red = 8'hcc;    Green = 8'hc2;    Blue = 8'h66;
end 13'h9b2:    begin Red = 8'ha1;    Green = 8'hac;    Blue = 8'h4c;
end 13'h9b3:    begin Red = 8'h63;    Green = 8'h58;    Blue = 8'h57;
end 13'h9b4:    begin Red = 8'h80;    Green = 8'ha7;    Blue = 8'h42;
end 13'h9b5:    begin Red = 8'h7d;    Green = 8'h9d;    Blue = 8'h6d;
end 13'h9b6:    begin Red = 8'h88;    Green = 8'hb7;    Blue = 8'h8f;
end 13'h9b7:    begin Red = 8'h8a;    Green = 8'haf;    Blue = 8'h7c;
end 13'h9b8:    begin Red = 8'ha4;    Green = 8'h85;    Blue = 8'h51;
end 13'h9b9:    begin Red = 8'h75;    Green = 8'h71;    Blue = 8'h45;
end 13'h9ba:    begin Red = 8'h78;    Green = 8'h74;    Blue = 8'h57;
end 13'h9bb:    begin Red = 8'ha8;    Green = 8'h81;    Blue = 8'h5f;
end 13'h9bc:    begin Red = 8'h66;    Green = 8'h71;    Blue = 8'h5c;
end 13'h9bd:    begin Red = 8'h75;    Green = 8'h9b;    Blue = 8'h6f;
end 13'h9be:    begin Red = 8'h72;    Green = 8'ha5;    Blue = 8'h75;
end 13'h9bf:    begin Red = 8'h83;    Green = 8'h6f;    Blue = 8'h4e;
end 13'h9c0:    begin Red = 8'h6d;    Green = 8'h6c;    Blue = 8'h3d;
end 13'h9c1:    begin Red = 8'hd6;    Green = 8'hc7;    Blue = 8'hac;
end 13'h9c2:    begin Red = 8'h8c;    Green = 8'h92;    Blue = 8'h73;
end 13'h9c3:    begin Red = 8'h7b;    Green = 8'h7f;    Blue = 8'h6c;
end 13'h9c4:    begin Red = 8'hc7;    Green = 8'hc1;    Blue = 8'ha2;
end 13'h9c5:    begin Red = 8'hde;    Green = 8'hc7;    Blue = 8'ha1;
end 13'h9c6:    begin Red = 8'hd7;    Green = 8'hbe;    Blue = 8'h9a;
end 13'h9c7:    begin Red = 8'he7;    Green = 8'hd2;    Blue = 8'hae;
end 13'h9c8:    begin Red = 8'hd2;    Green = 8'hb8;    Blue = 8'h96;
end 13'h9c9:    begin Red = 8'hae;    Green = 8'h9e;    Blue = 8'h76;
end 13'h9ca:    begin Red = 8'hff;    Green = 8'hf8;    Blue = 8'hdc;
end 13'h9cb:    begin Red = 8'hd6;    Green = 8'hc3;    Blue = 8'h95;
end 13'h9cc:    begin Red = 8'h6c;    Green = 8'h75;    Blue = 8'h5d;
end 13'h9cd:    begin Red = 8'hac;    Green = 8'h87;    Blue = 8'h51;
end 13'h9ce:    begin Red = 8'h71;    Green = 8'h75;    Blue = 8'h5d;
end 13'h9cf:    begin Red = 8'h98;    Green = 8'h70;    Blue = 8'h46;
end 13'h9d0:    begin Red = 8'hf5;    Green = 8'hda;    Blue = 8'hb7;
end 13'h9d1:    begin Red = 8'hd7;    Green = 8'hc2;    Blue = 8'h9e;
end 13'h9d2:    begin Red = 8'hbe;    Green = 8'hc4;    Blue = 8'hb6;
end 13'h9d3:    begin Red = 8'hb2;    Green = 8'hc4;    Blue = 8'hbf;
end 13'h9d4:    begin Red = 8'hcc;    Green = 8'hde;    Blue = 8'hd9;
end 13'h9d5:    begin Red = 8'h93;    Green = 8'h8d;    Blue = 8'h7e;
end 13'h9d6:    begin Red = 8'h90;    Green = 8'h8b;    Blue = 8'h7c;
end 13'h9d7:    begin Red = 8'h98;    Green = 8'h94;    Blue = 8'h82;
end 13'h9d8:    begin Red = 8'h9b;    Green = 8'h95;    Blue = 8'h84;
end 13'h9d9:    begin Red = 8'ha0;    Green = 8'h9a;    Blue = 8'h89;
end 13'h9da:    begin Red = 8'hca;    Green = 8'hcb;    Blue = 8'h49;
end 13'h9db:    begin Red = 8'h5d;    Green = 8'h69;    Blue = 8'h51;
end 13'h9dc:    begin Red = 8'hd8;    Green = 8'hd4;    Blue = 8'h5a;
end 13'h9dd:    begin Red = 8'hd3;    Green = 8'hd0;    Blue = 8'h65;
end 13'h9de:    begin Red = 8'hb9;    Green = 8'hd6;    Blue = 8'h49;
end 13'h9df:    begin Red = 8'h5e;    Green = 8'h4e;    Blue = 8'h5b;
end 13'h9e0:    begin Red = 8'h68;    Green = 8'h5f;    Blue = 8'h5a;
end 13'h9e1:    begin Red = 8'had;    Green = 8'hc7;    Blue = 8'h40;
end 13'h9e2:    begin Red = 8'ha2;    Green = 8'h6e;    Blue = 8'h5d;
end 13'h9e3:    begin Red = 8'hae;    Green = 8'h86;    Blue = 8'h5f;
end 13'h9e4:    begin Red = 8'hb8;    Green = 8'h88;    Blue = 8'h5a;
end 13'h9e5:    begin Red = 8'h62;    Green = 8'h73;    Blue = 8'h59;
end 13'h9e6:    begin Red = 8'h65;    Green = 8'h71;    Blue = 8'h61;
end 13'h9e7:    begin Red = 8'h64;    Green = 8'h6a;    Blue = 8'h5a;
end 13'h9e8:    begin Red = 8'ha1;    Green = 8'h76;    Blue = 8'h53;
end 13'h9e9:    begin Red = 8'hdf;    Green = 8'hbb;    Blue = 8'h93;
end 13'h9ea:    begin Red = 8'hc1;    Green = 8'hbd;    Blue = 8'h9d;
end 13'h9eb:    begin Red = 8'h81;    Green = 8'h86;    Blue = 8'h6b;
end 13'h9ec:    begin Red = 8'hce;    Green = 8'hb7;    Blue = 8'h90;
end 13'h9ed:    begin Red = 8'he7;    Green = 8'hd0;    Blue = 8'hb8;
end 13'h9ee:    begin Red = 8'hff;    Green = 8'hf0;    Blue = 8'hc3;
end 13'h9ef:    begin Red = 8'ha7;    Green = 8'h87;    Blue = 8'h5d;
end 13'h9f0:    begin Red = 8'h79;    Green = 8'h75;    Blue = 8'h46;
end 13'h9f1:    begin Red = 8'hb3;    Green = 8'h86;    Blue = 8'h55;
end 13'h9f2:    begin Red = 8'h62;    Green = 8'h72;    Blue = 8'h5d;
end 13'h9f3:    begin Red = 8'h95;    Green = 8'h78;    Blue = 8'h52;
end 13'h9f4:    begin Red = 8'h9d;    Green = 8'h75;    Blue = 8'h58;
end 13'h9f5:    begin Red = 8'hed;    Green = 8'hda;    Blue = 8'hc2;
end 13'h9f6:    begin Red = 8'he4;    Green = 8'hcd;    Blue = 8'hb2;
end 13'h9f7:    begin Red = 8'hbf;    Green = 8'hb4;    Blue = 8'hbe;
end 13'h9f8:    begin Red = 8'h8a;    Green = 8'h83;    Blue = 8'h75;
end 13'h9f9:    begin Red = 8'h91;    Green = 8'h8b;    Blue = 8'h78;
end 13'h9fa:    begin Red = 8'h94;    Green = 8'h90;    Blue = 8'h7d;
end 13'h9fb:    begin Red = 8'h98;    Green = 8'h93;    Blue = 8'h7e;
end 13'h9fc:    begin Red = 8'hcf;    Green = 8'hbe;    Blue = 8'h4a;
end 13'h9fd:    begin Red = 8'hc8;    Green = 8'hbb;    Blue = 8'h53;
end 13'h9fe:    begin Red = 8'ha4;    Green = 8'hbf;    Blue = 8'h51;
end 13'h9ff:    begin Red = 8'h8f;    Green = 8'h83;    Blue = 8'h4f;
end 13'ha00:    begin Red = 8'hb2;    Green = 8'h85;    Blue = 8'h60;
end 13'ha01:    begin Red = 8'h76;    Green = 8'h80;    Blue = 8'h69;
end 13'ha02:    begin Red = 8'h7a;    Green = 8'h7b;    Blue = 8'h6c;
end 13'ha03:    begin Red = 8'ha0;    Green = 8'h7e;    Blue = 8'h56;
end 13'ha04:    begin Red = 8'h69;    Green = 8'h73;    Blue = 8'h60;
end 13'ha05:    begin Red = 8'h6f;    Green = 8'h76;    Blue = 8'h5f;
end 13'ha06:    begin Red = 8'h6c;    Green = 8'h72;    Blue = 8'h65;
end 13'ha07:    begin Red = 8'h78;    Green = 8'h78;    Blue = 8'h6c;
end 13'ha08:    begin Red = 8'h79;    Green = 8'h75;    Blue = 8'h4b;
end 13'ha09:    begin Red = 8'h6e;    Green = 8'h71;    Blue = 8'h5f;
end 13'ha0a:    begin Red = 8'hd2;    Green = 8'hc0;    Blue = 8'h9f;
end 13'ha0b:    begin Red = 8'hd3;    Green = 8'hb6;    Blue = 8'h9f;
end 13'ha0c:    begin Red = 8'hd4;    Green = 8'hbd;    Blue = 8'ha2;
end 13'ha0d:    begin Red = 8'hd0;    Green = 8'hc0;    Blue = 8'ha4;
end 13'ha0e:    begin Red = 8'hc6;    Green = 8'hb4;    Blue = 8'h87;
end 13'ha0f:    begin Red = 8'ha3;    Green = 8'h8c;    Blue = 8'h71;
end 13'ha10:    begin Red = 8'he0;    Green = 8'hc6;    Blue = 8'ha3;
end 13'ha11:    begin Red = 8'h8f;    Green = 8'h79;    Blue = 8'h44;
end 13'ha12:    begin Red = 8'h64;    Green = 8'h75;    Blue = 8'h5c;
end 13'ha13:    begin Red = 8'h72;    Green = 8'h75;    Blue = 8'h67;
end 13'ha14:    begin Red = 8'h9e;    Green = 8'h90;    Blue = 8'h6d;
end 13'ha15:    begin Red = 8'h93;    Green = 8'h72;    Blue = 8'h4e;
end 13'ha16:    begin Red = 8'h9b;    Green = 8'h7b;    Blue = 8'h52;
end 13'ha17:    begin Red = 8'hca;    Green = 8'hb5;    Blue = 8'h8b;
end 13'ha18:    begin Red = 8'hd5;    Green = 8'hc8;    Blue = 8'ha1;
end 13'ha19:    begin Red = 8'hd6;    Green = 8'hbb;    Blue = 8'h9b;
end 13'ha1a:    begin Red = 8'hb8;    Green = 8'hbe;    Blue = 8'hc7;
end 13'ha1b:    begin Red = 8'hcf;    Green = 8'h91;    Blue = 8'hc1;
end 13'ha1c:    begin Red = 8'haf;    Green = 8'ha9;    Blue = 8'h9a;
end 13'ha1d:    begin Red = 8'hb3;    Green = 8'haf;    Blue = 8'h9d;
end 13'ha1e:    begin Red = 8'hb9;    Green = 8'hb3;    Blue = 8'ha2;
end 13'ha1f:    begin Red = 8'h9a;    Green = 8'h95;    Blue = 8'h80;
end 13'ha20:    begin Red = 8'hc7;    Green = 8'hb7;    Blue = 8'h5d;
end 13'ha21:    begin Red = 8'h59;    Green = 8'h4e;    Blue = 8'h3f;
end 13'ha22:    begin Red = 8'h65;    Green = 8'h65;    Blue = 8'h4c;
end 13'ha23:    begin Red = 8'h57;    Green = 8'h63;    Blue = 8'h49;
end 13'ha24:    begin Red = 8'hec;    Green = 8'hc5;    Blue = 8'ha3;
end 13'ha25:    begin Red = 8'he8;    Green = 8'hb7;    Blue = 8'h94;
end 13'ha26:    begin Red = 8'h7a;    Green = 8'h72;    Blue = 8'h5e;
end 13'ha27:    begin Red = 8'h91;    Green = 8'h75;    Blue = 8'h64;
end 13'ha28:    begin Red = 8'h7c;    Green = 8'h75;    Blue = 8'h3f;
end 13'ha29:    begin Red = 8'h8d;    Green = 8'h76;    Blue = 8'h48;
end 13'ha2a:    begin Red = 8'h6d;    Green = 8'h68;    Blue = 8'h3f;
end 13'ha2b:    begin Red = 8'haf;    Green = 8'hb7;    Blue = 8'h94;
end 13'ha2c:    begin Red = 8'h88;    Green = 8'h8b;    Blue = 8'h77;
end 13'ha2d:    begin Red = 8'h8e;    Green = 8'h92;    Blue = 8'h78;
end 13'ha2e:    begin Red = 8'he5;    Green = 8'hd4;    Blue = 8'had;
end 13'ha2f:    begin Red = 8'h52;    Green = 8'h47;    Blue = 8'h47;
end 13'ha30:    begin Red = 8'h52;    Green = 8'h4a;    Blue = 8'h4d;
end 13'ha31:    begin Red = 8'h4f;    Green = 8'h49;    Blue = 8'h47;
end 13'ha32:    begin Red = 8'h98;    Green = 8'h87;    Blue = 8'h68;
end 13'ha33:    begin Red = 8'h58;    Green = 8'h4d;    Blue = 8'h4d;
end 13'ha34:    begin Red = 8'h55;    Green = 8'h4a;    Blue = 8'h4a;
end 13'ha35:    begin Red = 8'h41;    Green = 8'h35;    Blue = 8'h37;
end 13'ha36:    begin Red = 8'hf6;    Green = 8'he1;    Blue = 8'hba;
end 13'ha37:    begin Red = 8'h51;    Green = 8'h48;    Blue = 8'h4b;
end 13'ha38:    begin Red = 8'h55;    Green = 8'h47;    Blue = 8'h4c;
end 13'ha39:    begin Red = 8'h5b;    Green = 8'h46;    Blue = 8'h4e;
end 13'ha3a:    begin Red = 8'h9b;    Green = 8'hb3;    Blue = 8'h8a;
end 13'ha3b:    begin Red = 8'h9c;    Green = 8'ha5;    Blue = 8'h83;
end 13'ha3c:    begin Red = 8'h98;    Green = 8'ha0;    Blue = 8'h7e;
end 13'ha3d:    begin Red = 8'h98;    Green = 8'h9c;    Blue = 8'h79;
end 13'ha3e:    begin Red = 8'hfd;    Green = 8'hf4;    Blue = 8'hcf;
end 13'ha3f:    begin Red = 8'h51;    Green = 8'h3f;    Blue = 8'h4a;
end 13'ha40:    begin Red = 8'he5;    Green = 8'hd2;    Blue = 8'hb1;
end 13'ha41:    begin Red = 8'hc2;    Green = 8'hbc;    Blue = 8'hc3;
end 13'ha42:    begin Red = 8'hc7;    Green = 8'h86;    Blue = 8'hb9;
end 13'ha43:    begin Red = 8'haa;    Green = 8'ha5;    Blue = 8'h92;
end 13'ha44:    begin Red = 8'hac;    Green = 8'ha7;    Blue = 8'h94;
end 13'ha45:    begin Red = 8'h84;    Green = 8'h7f;    Blue = 8'h70;
end 13'ha46:    begin Red = 8'h83;    Green = 8'h7e;    Blue = 8'h6c;
end 13'ha47:    begin Red = 8'h87;    Green = 8'h81;    Blue = 8'h73;
end 13'ha48:    begin Red = 8'h78;    Green = 8'h83;    Blue = 8'h3d;
end 13'ha49:    begin Red = 8'h83;    Green = 8'h88;    Blue = 8'h4d;
end 13'ha4a:    begin Red = 8'h67;    Green = 8'h70;    Blue = 8'h50;
end 13'ha4b:    begin Red = 8'h4f;    Green = 8'h61;    Blue = 8'h3d;
end 13'ha4c:    begin Red = 8'h63;    Green = 8'h71;    Blue = 8'h46;
end 13'ha4d:    begin Red = 8'hd0;    Green = 8'ha0;    Blue = 8'h7a;
end 13'ha4e:    begin Red = 8'hcb;    Green = 8'h9b;    Blue = 8'h74;
end 13'ha4f:    begin Red = 8'h8c;    Green = 8'h81;    Blue = 8'h64;
end 13'ha50:    begin Red = 8'hca;    Green = 8'h99;    Blue = 8'h71;
end 13'ha51:    begin Red = 8'h80;    Green = 8'h97;    Blue = 8'h51;
end 13'ha52:    begin Red = 8'hb3;    Green = 8'h88;    Blue = 8'h6c;
end 13'ha53:    begin Red = 8'h3e;    Green = 8'h38;    Blue = 8'h3f;
end 13'ha54:    begin Red = 8'h44;    Green = 8'h3c;    Blue = 8'h3b;
end 13'ha55:    begin Red = 8'h44;    Green = 8'h3c;    Blue = 8'h34;
end 13'ha56:    begin Red = 8'h46;    Green = 8'h42;    Blue = 8'h3f;
end 13'ha57:    begin Red = 8'h91;    Green = 8'h87;    Blue = 8'h6d;
end 13'ha58:    begin Red = 8'hed;    Green = 8'hb8;    Blue = 8'h96;
end 13'ha59:    begin Red = 8'h9b;    Green = 8'haf;    Blue = 8'h8e;
end 13'ha5a:    begin Red = 8'h66;    Green = 8'h6c;    Blue = 8'h4f;
end 13'ha5b:    begin Red = 8'h8b;    Green = 8'h7e;    Blue = 8'h6a;
end 13'ha5c:    begin Red = 8'h41;    Green = 8'h3d;    Blue = 8'h42;
end 13'ha5d:    begin Red = 8'h3a;    Green = 8'h40;    Blue = 8'h42;
end 13'ha5e:    begin Red = 8'h9c;    Green = 8'h78;    Blue = 8'h46;
end 13'ha5f:    begin Red = 8'h8f;    Green = 8'h85;    Blue = 8'h78;
end 13'ha60:    begin Red = 8'hbf;    Green = 8'ha0;    Blue = 8'h83;
end 13'ha61:    begin Red = 8'hbe;    Green = 8'ha2;    Blue = 8'h8c;
end 13'ha62:    begin Red = 8'he4;    Green = 8'hbd;    Blue = 8'h9c;
end 13'ha63:    begin Red = 8'ha8;    Green = 8'haf;    Blue = 8'h8c;
end 13'ha64:    begin Red = 8'h88;    Green = 8'h8b;    Blue = 8'h72;
end 13'ha65:    begin Red = 8'h6a;    Green = 8'h5c;    Blue = 8'h59;
end 13'ha66:    begin Red = 8'h68;    Green = 8'h5a;    Blue = 8'h58;
end 13'ha67:    begin Red = 8'hed;    Green = 8'hd8;    Blue = 8'hac;
end 13'ha68:    begin Red = 8'h6f;    Green = 8'h61;    Blue = 8'h5d;
end 13'ha69:    begin Red = 8'h69;    Green = 8'h5e;    Blue = 8'h57;
end 13'ha6a:    begin Red = 8'h70;    Green = 8'h60;    Blue = 8'h61;
end 13'ha6b:    begin Red = 8'h71;    Green = 8'h65;    Blue = 8'h5f;
end 13'ha6c:    begin Red = 8'ha9;    Green = 8'hb2;    Blue = 8'h84;
end 13'ha6d:    begin Red = 8'h9d;    Green = 8'ha3;    Blue = 8'h80;
end 13'ha6e:    begin Red = 8'h94;    Green = 8'h99;    Blue = 8'h7b;
end 13'ha6f:    begin Red = 8'h69;    Green = 8'h6c;    Blue = 8'h59;
end 13'ha70:    begin Red = 8'h97;    Green = 8'h75;    Blue = 8'h4a;
end 13'ha71:    begin Red = 8'hee;    Green = 8'hd7;    Blue = 8'ha7;
end 13'ha72:    begin Red = 8'h9c;    Green = 8'h86;    Blue = 8'h67;
end 13'ha73:    begin Red = 8'ha2;    Green = 8'h9c;    Blue = 8'h8e;
end 13'ha74:    begin Red = 8'ha7;    Green = 8'ha3;    Blue = 8'h90;
end 13'ha75:    begin Red = 8'hb0;    Green = 8'hac;    Blue = 8'h97;
end 13'ha76:    begin Red = 8'hb2;    Green = 8'had;    Blue = 8'h9b;
end 13'ha77:    begin Red = 8'h6c;    Green = 8'h7c;    Blue = 8'h55;
end 13'ha78:    begin Red = 8'h80;    Green = 8'h8a;    Blue = 8'h4e;
end 13'ha79:    begin Red = 8'h8b;    Green = 8'h75;    Blue = 8'h50;
end 13'ha7a:    begin Red = 8'h56;    Green = 8'h68;    Blue = 8'h43;
end 13'ha7b:    begin Red = 8'h5b;    Green = 8'h66;    Blue = 8'h4a;
end 13'ha7c:    begin Red = 8'h96;    Green = 8'h78;    Blue = 8'h57;
end 13'ha7d:    begin Red = 8'h4f;    Green = 8'h46;    Blue = 8'h42;
end 13'ha7e:    begin Red = 8'h92;    Green = 8'h80;    Blue = 8'h6d;
end 13'ha7f:    begin Red = 8'he7;    Green = 8'hb6;    Blue = 8'h90;
end 13'ha80:    begin Red = 8'h6a;    Green = 8'h6e;    Blue = 8'h55;
end 13'ha81:    begin Red = 8'hb5;    Green = 8'h9f;    Blue = 8'h81;
end 13'ha82:    begin Red = 8'had;    Green = 8'h9d;    Blue = 8'h81;
end 13'ha83:    begin Red = 8'hbb;    Green = 8'ha7;    Blue = 8'h80;
end 13'ha84:    begin Red = 8'h82;    Green = 8'h7c;    Blue = 8'h73;
end 13'ha85:    begin Red = 8'h9e;    Green = 8'h94;    Blue = 8'h86;
end 13'ha86:    begin Red = 8'h9d;    Green = 8'h94;    Blue = 8'h8a;
end 13'ha87:    begin Red = 8'h8c;    Green = 8'h7e;    Blue = 8'h76;
end 13'ha88:    begin Red = 8'h8a;    Green = 8'h80;    Blue = 8'h72;
end 13'ha89:    begin Red = 8'hab;    Green = 8'h9e;    Blue = 8'h92;
end 13'ha8a:    begin Red = 8'haa;    Green = 8'ha0;    Blue = 8'h90;
end 13'ha8b:    begin Red = 8'h97;    Green = 8'h8c;    Blue = 8'h86;
end 13'ha8c:    begin Red = 8'ha0;    Green = 8'h96;    Blue = 8'h88;
end 13'ha8d:    begin Red = 8'h9f;    Green = 8'h9a;    Blue = 8'h85;
end 13'ha8e:    begin Red = 8'had;    Green = 8'ha0;    Blue = 8'h96;
end 13'ha8f:    begin Red = 8'h9d;    Green = 8'haa;    Blue = 8'h78;
end 13'ha90:    begin Red = 8'ha5;    Green = 8'hac;    Blue = 8'h7f;
end 13'ha91:    begin Red = 8'hfc;    Green = 8'hf2;    Blue = 8'hd4;
end 13'ha92:    begin Red = 8'h92;    Green = 8'h87;    Blue = 8'h71;
end 13'ha93:    begin Red = 8'hbf;    Green = 8'hac;    Blue = 8'h7f;
end 13'ha94:    begin Red = 8'h9f;    Green = 8'h95;    Blue = 8'h82;
end 13'ha95:    begin Red = 8'hbf;    Green = 8'hc7;    Blue = 8'hcc;
end 13'ha96:    begin Red = 8'hd1;    Green = 8'hc5;    Blue = 8'h98;
end 13'ha97:    begin Red = 8'hd7;    Green = 8'hcb;    Blue = 8'h9e;
end 13'ha98:    begin Red = 8'hdc;    Green = 8'hd0;    Blue = 8'ha1;
end 13'ha99:    begin Red = 8'hda;    Green = 8'hcf;    Blue = 8'h9f;
end 13'ha9a:    begin Red = 8'hc4;    Green = 8'hbf;    Blue = 8'hab;
end 13'ha9b:    begin Red = 8'hc7;    Green = 8'hc3;    Blue = 8'hac;
end 13'ha9c:    begin Red = 8'hd2;    Green = 8'hce;    Blue = 8'hb7;
end 13'ha9d:    begin Red = 8'hd0;    Green = 8'hcc;    Blue = 8'hb5;
end 13'ha9e:    begin Red = 8'h92;    Green = 8'h8e;    Blue = 8'h76;
end 13'ha9f:    begin Red = 8'h65;    Green = 8'h6b;    Blue = 8'h44;
end 13'haa0:    begin Red = 8'h63;    Green = 8'h6c;    Blue = 8'h4d;
end 13'haa1:    begin Red = 8'h7b;    Green = 8'h88;    Blue = 8'h41;
end 13'haa2:    begin Red = 8'h76;    Green = 8'h8b;    Blue = 8'h52;
end 13'haa3:    begin Red = 8'h46;    Green = 8'h51;    Blue = 8'h39;
end 13'haa4:    begin Red = 8'hc6;    Green = 8'ha0;    Blue = 8'h78;
end 13'haa5:    begin Red = 8'hc5;    Green = 8'h96;    Blue = 8'h75;
end 13'haa6:    begin Red = 8'h82;    Green = 8'h7c;    Blue = 8'h5d;
end 13'haa7:    begin Red = 8'hc1;    Green = 8'h93;    Blue = 8'h6b;
end 13'haa8:    begin Red = 8'h74;    Green = 8'h7b;    Blue = 8'h4f;
end 13'haa9:    begin Red = 8'hbb;    Green = 8'h94;    Blue = 8'h6c;
end 13'haaa:    begin Red = 8'h5b;    Green = 8'h70;    Blue = 8'h37;
end 13'haab:    begin Red = 8'ha7;    Green = 8'h89;    Blue = 8'h64;
end 13'haac:    begin Red = 8'h8e;    Green = 8'h82;    Blue = 8'h6b;
end 13'haad:    begin Red = 8'ha3;    Green = 8'haa;    Blue = 8'h80;
end 13'haae:    begin Red = 8'hae;    Green = 8'hb5;    Blue = 8'h8b;
end 13'haaf:    begin Red = 8'h6d;    Green = 8'h5f;    Blue = 8'h55;
end 13'hab0:    begin Red = 8'hf0;    Green = 8'hce;    Blue = 8'haf;
end 13'hab1:    begin Red = 8'hab;    Green = 8'h9c;    Blue = 8'h7e;
end 13'hab2:    begin Red = 8'h7a;    Green = 8'h72;    Blue = 8'h6b;
end 13'hab3:    begin Red = 8'hb4;    Green = 8'ha2;    Blue = 8'h80;
end 13'hab4:    begin Red = 8'haa;    Green = 8'h9b;    Blue = 8'h81;
end 13'hab5:    begin Red = 8'h94;    Green = 8'h8a;    Blue = 8'h7d;
end 13'hab6:    begin Red = 8'h90;    Green = 8'h86;    Blue = 8'h73;
end 13'hab7:    begin Red = 8'ha8;    Green = 8'h99;    Blue = 8'h80;
end 13'hab8:    begin Red = 8'h9d;    Green = 8'ha7;    Blue = 8'h70;
end 13'hab9:    begin Red = 8'h9b;    Green = 8'ha1;    Blue = 8'h7a;
end 13'haba:    begin Red = 8'hf1;    Green = 8'he2;    Blue = 8'hc3;
end 13'habb:    begin Red = 8'h7f;    Green = 8'h7a;    Blue = 8'h65;
end 13'habc:    begin Red = 8'h9c;    Green = 8'h90;    Blue = 8'h79;
end 13'habd:    begin Red = 8'hae;    Green = 8'ha9;    Blue = 8'h96;
end 13'habe:    begin Red = 8'hb0;    Green = 8'hac;    Blue = 8'h9f;
end 13'habf:    begin Red = 8'hd5;    Green = 8'hc9;    Blue = 8'h9b;
end 13'hac0:    begin Red = 8'hd3;    Green = 8'hc7;    Blue = 8'h9d;
end 13'hac1:    begin Red = 8'hca;    Green = 8'hc1;    Blue = 8'h96;
end 13'hac2:    begin Red = 8'hd9;    Green = 8'hce;    Blue = 8'ha3;
end 13'hac3:    begin Red = 8'hde;    Green = 8'hd2;    Blue = 8'ha3;
end 13'hac4:    begin Red = 8'hc0;    Green = 8'hbb;    Blue = 8'ha7;
end 13'hac5:    begin Red = 8'hc4;    Green = 8'hbe;    Blue = 8'ha7;
end 13'hac6:    begin Red = 8'ha5;    Green = 8'hc3;    Blue = 8'ha6;
end 13'hac7:    begin Red = 8'h75;    Green = 8'h82;    Blue = 8'h56;
end 13'hac8:    begin Red = 8'h75;    Green = 8'h85;    Blue = 8'h58;
end 13'hac9:    begin Red = 8'h6d;    Green = 8'h80;    Blue = 8'h57;
end 13'haca:    begin Red = 8'h90;    Green = 8'h8b;    Blue = 8'h5d;
end 13'hacb:    begin Red = 8'h88;    Green = 8'h89;    Blue = 8'h53;
end 13'hacc:    begin Red = 8'h58;    Green = 8'h52;    Blue = 8'h44;
end 13'hacd:    begin Red = 8'hc3;    Green = 8'h99;    Blue = 8'h73;
end 13'hace:    begin Red = 8'h7d;    Green = 8'h7a;    Blue = 8'h55;
end 13'hacf:    begin Red = 8'h8e;    Green = 8'h86;    Blue = 8'h5f;
end 13'had0:    begin Red = 8'h84;    Green = 8'h83;    Blue = 8'h5a;
end 13'had1:    begin Red = 8'hc1;    Green = 8'h94;    Blue = 8'h70;
end 13'had2:    begin Red = 8'h93;    Green = 8'h85;    Blue = 8'h61;
end 13'had3:    begin Red = 8'hc1;    Green = 8'h9d;    Blue = 8'h71;
end 13'had4:    begin Red = 8'h65;    Green = 8'h5a;    Blue = 8'h42;
end 13'had5:    begin Red = 8'h60;    Green = 8'h58;    Blue = 8'h42;
end 13'had6:    begin Red = 8'h89;    Green = 8'ha7;    Blue = 8'h98;
end 13'had7:    begin Red = 8'h6b;    Green = 8'h78;    Blue = 8'h3f;
end 13'had8:    begin Red = 8'hac;    Green = 8'h88;    Blue = 8'h61;
end 13'had9:    begin Red = 8'h83;    Green = 8'h62;    Blue = 8'h51;
end 13'hada:    begin Red = 8'h7c;    Green = 8'h65;    Blue = 8'h5a;
end 13'hadb:    begin Red = 8'h92;    Green = 8'h81;    Blue = 8'h71;
end 13'hadc:    begin Red = 8'ha8;    Green = 8'hb0;    Blue = 8'h80;
end 13'hadd:    begin Red = 8'h84;    Green = 8'h76;    Blue = 8'h65;
end 13'hade:    begin Red = 8'he0;    Green = 8'hda;    Blue = 8'haf;
end 13'hadf:    begin Red = 8'he5;    Green = 8'hdf;    Blue = 8'hb3;
end 13'hae0:    begin Red = 8'ha9;    Green = 8'hb3;    Blue = 8'h8e;
end 13'hae1:    begin Red = 8'hea;    Green = 8'hd0;    Blue = 8'ha7;
end 13'hae2:    begin Red = 8'h7f;    Green = 8'h74;    Blue = 8'h6b;
end 13'hae3:    begin Red = 8'h6a;    Green = 8'h76;    Blue = 8'h95;
end 13'hae4:    begin Red = 8'h66;    Green = 8'h78;    Blue = 8'h9f;
end 13'hae5:    begin Red = 8'h68;    Green = 8'h78;    Blue = 8'h9c;
end 13'hae6:    begin Red = 8'h6c;    Green = 8'h7b;    Blue = 8'h99;
end 13'hae7:    begin Red = 8'h8d;    Green = 8'haf;    Blue = 8'hee;
end 13'hae8:    begin Red = 8'h94;    Green = 8'h88;    Blue = 8'h80;
end 13'hae9:    begin Red = 8'h85;    Green = 8'h7b;    Blue = 8'h74;
end 13'haea:    begin Red = 8'h70;    Green = 8'h86;    Blue = 8'hac;
end 13'haeb:    begin Red = 8'h73;    Green = 8'h80;    Blue = 8'hac;
end 13'haec:    begin Red = 8'h72;    Green = 8'h84;    Blue = 8'hab;
end 13'haed:    begin Red = 8'ha7;    Green = 8'hbb;    Blue = 8'hf2;
end 13'haee:    begin Red = 8'ha6;    Green = 8'h8a;    Blue = 8'h6c;
end 13'haef:    begin Red = 8'h99;    Green = 8'hb8;    Blue = 8'hf7;
end 13'haf0:    begin Red = 8'h6e;    Green = 8'h80;    Blue = 8'ha5;
end 13'haf1:    begin Red = 8'h74;    Green = 8'h83;    Blue = 8'ha3;
end 13'haf2:    begin Red = 8'ha7;    Green = 8'hac;    Blue = 8'h6e;
end 13'haf3:    begin Red = 8'heb;    Green = 8'hce;    Blue = 8'ha5;
end 13'haf4:    begin Red = 8'h65;    Green = 8'h76;    Blue = 8'h98;
end 13'haf5:    begin Red = 8'h68;    Green = 8'h79;    Blue = 8'ha7;
end 13'haf6:    begin Red = 8'h69;    Green = 8'h7c;    Blue = 8'h9c;
end 13'haf7:    begin Red = 8'h8e;    Green = 8'ha6;    Blue = 8'hdf;
end 13'haf8:    begin Red = 8'hc7;    Green = 8'h84;    Blue = 8'haf;
end 13'haf9:    begin Red = 8'hb3;    Green = 8'haa;    Blue = 8'h9f;
end 13'hafa:    begin Red = 8'ha0;    Green = 8'h94;    Blue = 8'h8e;
end 13'hafb:    begin Red = 8'he4;    Green = 8'hd8;    Blue = 8'hbe;
end 13'hafc:    begin Red = 8'h98;    Green = 8'h89;    Blue = 8'h88;
end 13'hafd:    begin Red = 8'ha3;    Green = 8'h98;    Blue = 8'h90;
end 13'hafe:    begin Red = 8'hd9;    Green = 8'hcc;    Blue = 8'h9c;
end 13'haff:    begin Red = 8'h6c;    Green = 8'h81;    Blue = 8'h61;
end 13'hb00:    begin Red = 8'h6b;    Green = 8'h5a;    Blue = 8'h4a;
end 13'hb01:    begin Red = 8'h8a;    Green = 8'h7c;    Blue = 8'h5c;
end 13'hb02:    begin Red = 8'haf;    Green = 8'h8e;    Blue = 8'h68;
end 13'hb03:    begin Red = 8'h5d;    Green = 8'h55;    Blue = 8'h3b;
end 13'hb04:    begin Red = 8'ha3;    Green = 8'h80;    Blue = 8'h5e;
end 13'hb05:    begin Red = 8'h43;    Green = 8'h40;    Blue = 8'h41;
end 13'hb06:    begin Red = 8'h4b;    Green = 8'h49;    Blue = 8'h42;
end 13'hb07:    begin Red = 8'h5a;    Green = 8'h51;    Blue = 8'h4a;
end 13'hb08:    begin Red = 8'hdc;    Green = 8'hb9;    Blue = 8'h9a;
end 13'hb09:    begin Red = 8'hd2;    Green = 8'ha7;    Blue = 8'h81;
end 13'hb0a:    begin Red = 8'h88;    Green = 8'h8d;    Blue = 8'h6a;
end 13'hb0b:    begin Red = 8'he2;    Green = 8'hde;    Blue = 8'haf;
end 13'hb0c:    begin Red = 8'he9;    Green = 8'he2;    Blue = 8'hbb;
end 13'hb0d:    begin Red = 8'hdc;    Green = 8'he2;    Blue = 8'hc0;
end 13'hb0e:    begin Red = 8'h74;    Green = 8'h77;    Blue = 8'h63;
end 13'hb0f:    begin Red = 8'hee;    Green = 8'he9;    Blue = 8'hc6;
end 13'hb10:    begin Red = 8'hd4;    Green = 8'hce;    Blue = 8'ha8;
end 13'hb11:    begin Red = 8'hbf;    Green = 8'hbb;    Blue = 8'h94;
end 13'hb12:    begin Red = 8'hbc;    Green = 8'hb7;    Blue = 8'h9b;
end 13'hb13:    begin Red = 8'h94;    Green = 8'h87;    Blue = 8'h7b;
end 13'hb14:    begin Red = 8'h80;    Green = 8'h7b;    Blue = 8'h6e;
end 13'hb15:    begin Red = 8'ha8;    Green = 8'h9b;    Blue = 8'h84;
end 13'hb16:    begin Red = 8'ha5;    Green = 8'h9b;    Blue = 8'h79;
end 13'hb17:    begin Red = 8'h9b;    Green = 8'h91;    Blue = 8'h7d;
end 13'hb18:    begin Red = 8'h95;    Green = 8'h90;    Blue = 8'h88;
end 13'hb19:    begin Red = 8'h8c;    Green = 8'h8e;    Blue = 8'h7b;
end 13'hb1a:    begin Red = 8'ha3;    Green = 8'h8a;    Blue = 8'h74;
end 13'hb1b:    begin Red = 8'hae;    Green = 8'h97;    Blue = 8'h74;
end 13'hb1c:    begin Red = 8'h9c;    Green = 8'hae;    Blue = 8'h7a;
end 13'hb1d:    begin Red = 8'ha1;    Green = 8'ha7;    Blue = 8'h80;
end 13'hb1e:    begin Red = 8'h7d;    Green = 8'h80;    Blue = 8'h66;
end 13'hb1f:    begin Red = 8'h84;    Green = 8'h88;    Blue = 8'h6c;
end 13'hb20:    begin Red = 8'h84;    Green = 8'h77;    Blue = 8'h71;
end 13'hb21:    begin Red = 8'h9e;    Green = 8'h8d;    Blue = 8'h78;
end 13'hb22:    begin Red = 8'hc6;    Green = 8'h90;    Blue = 8'hc6;
end 13'hb23:    begin Red = 8'he2;    Green = 8'ha0;    Blue = 8'hd1;
end 13'hb24:    begin Red = 8'hd4;    Green = 8'h9b;    Blue = 8'hd2;
end 13'hb25:    begin Red = 8'hdc;    Green = 8'h9b;    Blue = 8'hce;
end 13'hb26:    begin Red = 8'hc3;    Green = 8'hba;    Blue = 8'h8d;
end 13'hb27:    begin Red = 8'hc7;    Green = 8'hbf;    Blue = 8'h90;
end 13'hb28:    begin Red = 8'he1;    Green = 8'hd6;    Blue = 8'hbe;
end 13'hb29:    begin Red = 8'hb4;    Green = 8'ha9;    Blue = 8'h92;
end 13'hb2a:    begin Red = 8'hbf;    Green = 8'hb6;    Blue = 8'h96;
end 13'hb2b:    begin Red = 8'ha0;    Green = 8'h90;    Blue = 8'h95;
end 13'hb2c:    begin Red = 8'ha3;    Green = 8'hc3;    Blue = 8'hb2;
end 13'hb2d:    begin Red = 8'h5f;    Green = 8'h6d;    Blue = 8'h4f;
end 13'hb2e:    begin Red = 8'h8f;    Green = 8'h7a;    Blue = 8'h51;
end 13'hb2f:    begin Red = 8'h59;    Green = 8'h55;    Blue = 8'h37;
end 13'hb30:    begin Red = 8'h89;    Green = 8'h83;    Blue = 8'h4f;
end 13'hb31:    begin Red = 8'h60;    Green = 8'h55;    Blue = 8'h46;
end 13'hb32:    begin Red = 8'hbe;    Green = 8'h94;    Blue = 8'h72;
end 13'hb33:    begin Red = 8'h92;    Green = 8'h86;    Blue = 8'h5a;
end 13'hb34:    begin Red = 8'h90;    Green = 8'h8b;    Blue = 8'h63;
end 13'hb35:    begin Red = 8'h7d;    Green = 8'h70;    Blue = 8'h43;
end 13'hb36:    begin Red = 8'h72;    Green = 8'h63;    Blue = 8'h35;
end 13'hb37:    begin Red = 8'he5;    Green = 8'hc2;    Blue = 8'ha3;
end 13'hb38:    begin Red = 8'h98;    Green = 8'h7d;    Blue = 8'h5d;
end 13'hb39:    begin Red = 8'hec;    Green = 8'hc8;    Blue = 8'ha7;
end 13'hb3a:    begin Red = 8'ha7;    Green = 8'haf;    Blue = 8'h7d;
end 13'hb3b:    begin Red = 8'he1;    Green = 8'hdc;    Blue = 8'hac;
end 13'hb3c:    begin Red = 8'hd1;    Green = 8'hd6;    Blue = 8'hb3;
end 13'hb3d:    begin Red = 8'he2;    Green = 8'hdb;    Blue = 8'hb7;
end 13'hb3e:    begin Red = 8'he5;    Green = 8'he0;    Blue = 8'hbd;
end 13'hb3f:    begin Red = 8'hcf;    Green = 8'hc9;    Blue = 8'ha4;
end 13'hb40:    begin Red = 8'hba;    Green = 8'hb3;    Blue = 8'h97;
end 13'hb41:    begin Red = 8'he8;    Green = 8'hcf;    Blue = 8'ha4;
end 13'hb42:    begin Red = 8'h7e;    Green = 8'h71;    Blue = 8'h6a;
end 13'hb43:    begin Red = 8'h91;    Green = 8'h88;    Blue = 8'h87;
end 13'hb44:    begin Red = 8'h99;    Green = 8'h86;    Blue = 8'h84;
end 13'hb45:    begin Red = 8'h99;    Green = 8'h88;    Blue = 8'h7d;
end 13'hb46:    begin Red = 8'h98;    Green = 8'h8a;    Blue = 8'h82;
end 13'hb47:    begin Red = 8'he4;    Green = 8'hcc;    Blue = 8'ha4;
end 13'hb48:    begin Red = 8'h8c;    Green = 8'h7d;    Blue = 8'h71;
end 13'hb49:    begin Red = 8'h9f;    Green = 8'h98;    Blue = 8'h80;
end 13'hb4a:    begin Red = 8'h9e;    Green = 8'h98;    Blue = 8'h8a;
end 13'hb4b:    begin Red = 8'ha4;    Green = 8'h97;    Blue = 8'h8a;
end 13'hb4c:    begin Red = 8'ha7;    Green = 8'h90;    Blue = 8'h84;
end 13'hb4d:    begin Red = 8'h89;    Green = 8'h84;    Blue = 8'h7b;
end 13'hb4e:    begin Red = 8'ha1;    Green = 8'h93;    Blue = 8'h89;
end 13'hb4f:    begin Red = 8'ha3;    Green = 8'h94;    Blue = 8'h8b;
end 13'hb50:    begin Red = 8'h99;    Green = 8'ha3;    Blue = 8'h7d;
end 13'hb51:    begin Red = 8'h80;    Green = 8'h75;    Blue = 8'h6e;
end 13'hb52:    begin Red = 8'h94;    Green = 8'h8a;    Blue = 8'h85;
end 13'hb53:    begin Red = 8'hdc;    Green = 8'ha7;    Blue = 8'hd1;
end 13'hb54:    begin Red = 8'hdb;    Green = 8'ha4;    Blue = 8'hcf;
end 13'hb55:    begin Red = 8'hd6;    Green = 8'ha5;    Blue = 8'hca;
end 13'hb56:    begin Red = 8'hc0;    Green = 8'hb6;    Blue = 8'h92;
end 13'hb57:    begin Red = 8'h9b;    Green = 8'h90;    Blue = 8'h89;
end 13'hb58:    begin Red = 8'hb4;    Green = 8'ha8;    Blue = 8'h8e;
end 13'hb59:    begin Red = 8'hba;    Green = 8'hb0;    Blue = 8'h8f;
end 13'hb5a:    begin Red = 8'h9b;    Green = 8'h8d;    Blue = 8'h8c;
end 13'hb5b:    begin Red = 8'hd6;    Green = 8'hcd;    Blue = 8'ha2;
end 13'hb5c:    begin Red = 8'h68;    Green = 8'h69;    Blue = 8'h42;
end 13'hb5d:    begin Red = 8'h9b;    Green = 8'hac;    Blue = 8'h59;
end 13'hb5e:    begin Red = 8'h93;    Green = 8'ha7;    Blue = 8'h56;
end 13'hb5f:    begin Red = 8'hac;    Green = 8'h7d;    Blue = 8'h57;
end 13'hb60:    begin Red = 8'ha3;    Green = 8'h81;    Blue = 8'h57;
end 13'hb61:    begin Red = 8'h84;    Green = 8'h7a;    Blue = 8'h52;
end 13'hb62:    begin Red = 8'h84;    Green = 8'h7d;    Blue = 8'h4a;
end 13'hb63:    begin Red = 8'hbb;    Green = 8'h94;    Blue = 8'h74;
end 13'hb64:    begin Red = 8'h65;    Green = 8'h5d;    Blue = 8'h38;
end 13'hb65:    begin Red = 8'h60;    Green = 8'h56;    Blue = 8'h4a;
end 13'hb66:    begin Red = 8'he4;    Green = 8'hb4;    Blue = 8'h8b;
end 13'hb67:    begin Red = 8'h9b;    Green = 8'ha5;    Blue = 8'h7f;
end 13'hb68:    begin Red = 8'hac;    Green = 8'h85;    Blue = 8'h65;
end 13'hb69:    begin Red = 8'ha3;    Green = 8'h85;    Blue = 8'h61;
end 13'hb6a:    begin Red = 8'hde;    Green = 8'hc6;    Blue = 8'ha9;
end 13'hb6b:    begin Red = 8'hf7;    Green = 8'hde;    Blue = 8'hb3;
end 13'hb6c:    begin Red = 8'h69;    Green = 8'h7a;    Blue = 8'ha0;
end 13'hb6d:    begin Red = 8'h65;    Green = 8'h7c;    Blue = 8'h94;
end 13'hb6e:    begin Red = 8'h98;    Green = 8'hb7;    Blue = 8'hf2;
end 13'hb6f:    begin Red = 8'h92;    Green = 8'ha8;    Blue = 8'he3;
end 13'hb70:    begin Red = 8'h92;    Green = 8'h84;    Blue = 8'h64;
end 13'hb71:    begin Red = 8'he2;    Green = 8'hca;    Blue = 8'haf;
end 13'hb72:    begin Red = 8'h72;    Green = 8'h83;    Blue = 8'ha7;
end 13'hb73:    begin Red = 8'h71;    Green = 8'h82;    Blue = 8'hb4;
end 13'hb74:    begin Red = 8'h70;    Green = 8'h84;    Blue = 8'ha4;
end 13'hb75:    begin Red = 8'h9e;    Green = 8'hbb;    Blue = 8'hf6;
end 13'hb76:    begin Red = 8'h96;    Green = 8'hbb;    Blue = 8'hf3;
end 13'hb77:    begin Red = 8'h9b;    Green = 8'hbf;    Blue = 8'hf5;
end 13'hb78:    begin Red = 8'h9f;    Green = 8'hbb;    Blue = 8'hfb;
end 13'hb79:    begin Red = 8'ha9;    Green = 8'hc8;    Blue = 8'hfd;
end 13'hb7a:    begin Red = 8'h72;    Green = 8'h88;    Blue = 8'had;
end 13'hb7b:    begin Red = 8'h78;    Green = 8'h83;    Blue = 8'haa;
end 13'hb7c:    begin Red = 8'h81;    Green = 8'h76;    Blue = 8'h74;
end 13'hb7d:    begin Red = 8'h6f;    Green = 8'h78;    Blue = 8'h9c;
end 13'hb7e:    begin Red = 8'h94;    Green = 8'hb3;    Blue = 8'hee;
end 13'hb7f:    begin Red = 8'h90;    Green = 8'ha7;    Blue = 8'he6;
end 13'hb80:    begin Red = 8'h90;    Green = 8'hab;    Blue = 8'he4;
end 13'hb81:    begin Red = 8'h91;    Green = 8'h88;    Blue = 8'h76;
end 13'hb82:    begin Red = 8'hb9;    Green = 8'hb9;    Blue = 8'hb9;
end 13'hb83:    begin Red = 8'h99;    Green = 8'h8e;    Blue = 8'h85;
end 13'hb84:    begin Red = 8'he7;    Green = 8'hdc;    Blue = 8'hc7;
end 13'hb85:    begin Red = 8'ha6;    Green = 8'h99;    Blue = 8'h8f;
end 13'hb86:    begin Red = 8'hc7;    Green = 8'hbe;    Blue = 8'ha9;
end 13'hb87:    begin Red = 8'h4d;    Green = 8'h4f;    Blue = 8'h42;
end 13'hb88:    begin Red = 8'h94;    Green = 8'ha4;    Blue = 8'h52;
end 13'hb89:    begin Red = 8'h41;    Green = 8'h44;    Blue = 8'h38;
end 13'hb8a:    begin Red = 8'h54;    Green = 8'h57;    Blue = 8'h43;
end 13'hb8b:    begin Red = 8'ha3;    Green = 8'hb9;    Blue = 8'h51;
end 13'hb8c:    begin Red = 8'hb0;    Green = 8'h8d;    Blue = 8'h5d;
end 13'hb8d:    begin Red = 8'h9b;    Green = 8'h78;    Blue = 8'h55;
end 13'hb8e:    begin Red = 8'h92;    Green = 8'h70;    Blue = 8'h47;
end 13'hb8f:    begin Red = 8'hd6;    Green = 8'hb7;    Blue = 8'h8c;
end 13'hb90:    begin Red = 8'h7e;    Green = 8'h8c;    Blue = 8'h6c;
end 13'hb91:    begin Red = 8'h93;    Green = 8'h99;    Blue = 8'h74;
end 13'hb92:    begin Red = 8'hed;    Green = 8'he7;    Blue = 8'hc3;
end 13'hb93:    begin Red = 8'hed;    Green = 8'he4;    Blue = 8'hc0;
end 13'hb94:    begin Red = 8'hbb;    Green = 8'hbe;    Blue = 8'ha0;
end 13'hb95:    begin Red = 8'hf0;    Green = 8'heb;    Blue = 8'hc5;
end 13'hb96:    begin Red = 8'hd8;    Green = 8'hd2;    Blue = 8'hac;
end 13'hb97:    begin Red = 8'h61;    Green = 8'h7c;    Blue = 8'h98;
end 13'hb98:    begin Red = 8'h6c;    Green = 8'h79;    Blue = 8'ha8;
end 13'hb99:    begin Red = 8'h94;    Green = 8'hb4;    Blue = 8'hf8;
end 13'hb9a:    begin Red = 8'h8c;    Green = 8'ha9;    Blue = 8'hef;
end 13'hb9b:    begin Red = 8'h94;    Green = 8'haa;    Blue = 8'hdf;
end 13'hb9c:    begin Red = 8'h8b;    Green = 8'h79;    Blue = 8'h6e;
end 13'hb9d:    begin Red = 8'h70;    Green = 8'h82;    Blue = 8'haa;
end 13'hb9e:    begin Red = 8'h74;    Green = 8'h85;    Blue = 8'ha6;
end 13'hb9f:    begin Red = 8'ha0;    Green = 8'h89;    Blue = 8'h6a;
end 13'hba0:    begin Red = 8'h93;    Green = 8'h86;    Blue = 8'h88;
end 13'hba1:    begin Red = 8'h9b;    Green = 8'hb8;    Blue = 8'hfe;
end 13'hba2:    begin Red = 8'h8c;    Green = 8'hac;    Blue = 8'he7;
end 13'hba3:    begin Red = 8'h88;    Green = 8'hab;    Blue = 8'he2;
end 13'hba4:    begin Red = 8'hc3;    Green = 8'hbe;    Blue = 8'hc6;
end 13'hba5:    begin Red = 8'hb5;    Green = 8'hbf;    Blue = 8'hb7;
end 13'hba6:    begin Red = 8'hc6;    Green = 8'hbe;    Blue = 8'h93;
end 13'hba7:    begin Red = 8'h91;    Green = 8'h87;    Blue = 8'h82;
end 13'hba8:    begin Red = 8'h96;    Green = 8'h89;    Blue = 8'h8c;
end 13'hba9:    begin Red = 8'hf6;    Green = 8'hed;    Blue = 8'hcd;
end 13'hbaa:    begin Red = 8'h9a;    Green = 8'hb6;    Blue = 8'ha6;
end 13'hbab:    begin Red = 8'h92;    Green = 8'ha7;    Blue = 8'h3f;
end 13'hbac:    begin Red = 8'h49;    Green = 8'h4e;    Blue = 8'h36;
end 13'hbad:    begin Red = 8'h3b;    Green = 8'h3a;    Blue = 8'h39;
end 13'hbae:    begin Red = 8'ha2;    Green = 8'hb8;    Blue = 8'h56;
end 13'hbaf:    begin Red = 8'hae;    Green = 8'hc6;    Blue = 8'h5e;
end 13'hbb0:    begin Red = 8'h90;    Green = 8'h7e;    Blue = 8'h50;
end 13'hbb1:    begin Red = 8'h89;    Green = 8'h7b;    Blue = 8'h53;
end 13'hbb2:    begin Red = 8'h80;    Green = 8'h75;    Blue = 8'h55;
end 13'hbb3:    begin Red = 8'h9f;    Green = 8'h81;    Blue = 8'h58;
end 13'hbb4:    begin Red = 8'haf;    Green = 8'h8b;    Blue = 8'h5b;
end 13'hbb5:    begin Red = 8'h5f;    Green = 8'h52;    Blue = 8'h38;
end 13'hbb6:    begin Red = 8'ha2;    Green = 8'h7c;    Blue = 8'h55;
end 13'hbb7:    begin Red = 8'h9d;    Green = 8'h74;    Blue = 8'h46;
end 13'hbb8:    begin Red = 8'h97;    Green = 8'h6b;    Blue = 8'h40;
end 13'hbb9:    begin Red = 8'h8d;    Green = 8'ha0;    Blue = 8'h76;
end 13'hbba:    begin Red = 8'haf;    Green = 8'hab;    Blue = 8'h91;
end 13'hbbb:    begin Red = 8'h9f;    Green = 8'ha2;    Blue = 8'h88;
end 13'hbbc:    begin Red = 8'ha8;    Green = 8'haa;    Blue = 8'h8c;
end 13'hbbd:    begin Red = 8'hb2;    Green = 8'had;    Blue = 8'h92;
end 13'hbbe:    begin Red = 8'h94;    Green = 8'h8f;    Blue = 8'h78;
end 13'hbbf:    begin Red = 8'h96;    Green = 8'hb4;    Blue = 8'hf5;
end 13'hbc0:    begin Red = 8'h85;    Green = 8'h7a;    Blue = 8'h70;
end 13'hbc1:    begin Red = 8'hf5;    Green = 8'hdd;    Blue = 8'hb5;
end 13'hbc2:    begin Red = 8'hbd;    Green = 8'hc5;    Blue = 8'hb2;
end 13'hbc3:    begin Red = 8'hd7;    Green = 8'ha8;    Blue = 8'hcd;
end 13'hbc4:    begin Red = 8'hca;    Green = 8'hba;    Blue = 8'h91;
end 13'hbc5:    begin Red = 8'h99;    Green = 8'hb4;    Blue = 8'ha1;
end 13'hbc6:    begin Red = 8'h65;    Green = 8'h70;    Blue = 8'h4b;
end 13'hbc7:    begin Red = 8'h5b;    Green = 8'h5b;    Blue = 8'h46;
end 13'hbc8:    begin Red = 8'h50;    Green = 8'h52;    Blue = 8'h43;
end 13'hbc9:    begin Red = 8'h69;    Green = 8'h6d;    Blue = 8'h49;
end 13'hbca:    begin Red = 8'h7a;    Green = 8'h72;    Blue = 8'h4a;
end 13'hbcb:    begin Red = 8'h73;    Green = 8'h96;    Blue = 8'h84;
end 13'hbcc:    begin Red = 8'had;    Green = 8'h9a;    Blue = 8'h75;
end 13'hbcd:    begin Red = 8'h49;    Green = 8'h47;    Blue = 8'h3e;
end 13'hbce:    begin Red = 8'h5b;    Green = 8'h55;    Blue = 8'h47;
end 13'hbcf:    begin Red = 8'h79;    Green = 8'h8c;    Blue = 8'h6a;
end 13'hbd0:    begin Red = 8'h74;    Green = 8'h79;    Blue = 8'h5f;
end 13'hbd1:    begin Red = 8'h84;    Green = 8'h73;    Blue = 8'h68;
end 13'hbd2:    begin Red = 8'h90;    Green = 8'h80;    Blue = 8'h6a;
end 13'hbd3:    begin Red = 8'h9f;    Green = 8'h90;    Blue = 8'h76;
end 13'hbd4:    begin Red = 8'he7;    Green = 8'he2;    Blue = 8'hb3;
end 13'hbd5:    begin Red = 8'hbd;    Green = 8'hc4;    Blue = 8'ha0;
end 13'hbd6:    begin Red = 8'h98;    Green = 8'h99;    Blue = 8'h80;
end 13'hbd7:    begin Red = 8'ha5;    Green = 8'h9e;    Blue = 8'h87;
end 13'hbd8:    begin Red = 8'hac;    Green = 8'hb3;    Blue = 8'h90;
end 13'hbd9:    begin Red = 8'h8a;    Green = 8'h8d;    Blue = 8'h73;
end 13'hbda:    begin Red = 8'hfd;    Green = 8'hf0;    Blue = 8'hcd;
end 13'hbdb:    begin Red = 8'hc1;    Green = 8'hb9;    Blue = 8'hc0;
end 13'hbdc:    begin Red = 8'hcb;    Green = 8'h8f;    Blue = 8'hb3;
end 13'hbdd:    begin Red = 8'hbc;    Green = 8'h84;    Blue = 8'hb6;
end 13'hbde:    begin Red = 8'hd3;    Green = 8'hcb;    Blue = 8'hd4;
end 13'hbdf:    begin Red = 8'hac;    Green = 8'hac;    Blue = 8'h99;
end 13'hbe0:    begin Red = 8'ha0;    Green = 8'h91;    Blue = 8'h90;
end 13'hbe1:    begin Red = 8'hde;    Green = 8'hd4;    Blue = 8'hb0;
end 13'hbe2:    begin Red = 8'hc6;    Green = 8'hb7;    Blue = 8'ha9;
end 13'hbe3:    begin Red = 8'h9b;    Green = 8'hc5;    Blue = 8'had;
end 13'hbe4:    begin Red = 8'h8a;    Green = 8'h88;    Blue = 8'h4b;
end 13'hbe5:    begin Red = 8'h82;    Green = 8'h80;    Blue = 8'h45;
end 13'hbe6:    begin Red = 8'h96;    Green = 8'haf;    Blue = 8'h6f;
end 13'hbe7:    begin Red = 8'h8b;    Green = 8'ha2;    Blue = 8'h5f;
end 13'hbe8:    begin Red = 8'h5b;    Green = 8'h5a;    Blue = 8'h4f;
end 13'hbe9:    begin Red = 8'h59;    Green = 8'h56;    Blue = 8'h4f;
end 13'hbea:    begin Red = 8'h65;    Green = 8'h77;    Blue = 8'h4c;
end 13'hbeb:    begin Red = 8'h71;    Green = 8'h7d;    Blue = 8'h43;
end 13'hbec:    begin Red = 8'h6d;    Green = 8'h75;    Blue = 8'h61;
end 13'hbed:    begin Red = 8'h81;    Green = 8'h6d;    Blue = 8'h39;
end 13'hbee:    begin Red = 8'h79;    Green = 8'h78;    Blue = 8'h49;
end 13'hbef:    begin Red = 8'ha3;    Green = 8'h77;    Blue = 8'h4e;
end 13'hbf0:    begin Red = 8'h93;    Green = 8'h6c;    Blue = 8'h46;
end 13'hbf1:    begin Red = 8'haf;    Green = 8'h86;    Blue = 8'h64;
end 13'hbf2:    begin Red = 8'h90;    Green = 8'h81;    Blue = 8'h74;
end 13'hbf3:    begin Red = 8'haf;    Green = 8'hb6;    Blue = 8'h90;
end 13'hbf4:    begin Red = 8'ha7;    Green = 8'h82;    Blue = 8'h5b;
end 13'hbf5:    begin Red = 8'h82;    Green = 8'h82;    Blue = 8'h6c;
end 13'hbf6:    begin Red = 8'hbe;    Green = 8'h86;    Blue = 8'hb8;
end 13'hbf7:    begin Red = 8'hce;    Green = 8'hd3;    Blue = 8'hd9;
end 13'hbf8:    begin Red = 8'hd6;    Green = 8'ha0;    Blue = 8'hc9;
end 13'hbf9:    begin Red = 8'hc1;    Green = 8'hbe;    Blue = 8'h93;
end 13'hbfa:    begin Red = 8'hc6;    Green = 8'hc1;    Blue = 8'h9b;
end 13'hbfb:    begin Red = 8'he0;    Green = 8'hd2;    Blue = 8'haa;
end 13'hbfc:    begin Red = 8'h84;    Green = 8'h80;    Blue = 8'h42;
end 13'hbfd:    begin Red = 8'h7a;    Green = 8'h73;    Blue = 8'h59;
end 13'hbfe:    begin Red = 8'h8c;    Green = 8'ha2;    Blue = 8'h65;
end 13'hbff:    begin Red = 8'h62;    Green = 8'h64;    Blue = 8'h51;
end 13'hc00:    begin Red = 8'h57;    Green = 8'h5a;    Blue = 8'h4d;
end 13'hc01:    begin Red = 8'h6f;    Green = 8'h80;    Blue = 8'h4c;
end 13'hc02:    begin Red = 8'h84;    Green = 8'h6d;    Blue = 8'h41;
end 13'hc03:    begin Red = 8'h80;    Green = 8'h6f;    Blue = 8'h51;
end 13'hc04:    begin Red = 8'h98;    Green = 8'h7d;    Blue = 8'h4a;
end 13'hc05:    begin Red = 8'hb2;    Green = 8'h92;    Blue = 8'h7d;
end 13'hc06:    begin Red = 8'had;    Green = 8'h95;    Blue = 8'h7a;
end 13'hc07:    begin Red = 8'hc7;    Green = 8'h90;    Blue = 8'hb9;
end 13'hc08:    begin Red = 8'hbf;    Green = 8'hb9;    Blue = 8'h9c;
end 13'hc09:    begin Red = 8'hce;    Green = 8'hc6;    Blue = 8'ha2;
end 13'hc0a:    begin Red = 8'h8f;    Green = 8'h90;    Blue = 8'h58;
end 13'hc0b:    begin Red = 8'h8a;    Green = 8'h85;    Blue = 8'h47;
end 13'hc0c:    begin Red = 8'h84;    Green = 8'h82;    Blue = 8'h47;
end 13'hc0d:    begin Red = 8'h71;    Green = 8'h70;    Blue = 8'h4d;
end 13'hc0e:    begin Red = 8'h75;    Green = 8'h84;    Blue = 8'h45;
end 13'hc0f:    begin Red = 8'h68;    Green = 8'h6e;    Blue = 8'h4e;
end 13'hc10:    begin Red = 8'h7a;    Green = 8'h8a;    Blue = 8'h45;
end 13'hc11:    begin Red = 8'h76;    Green = 8'h8d;    Blue = 8'h44;
end 13'hc12:    begin Red = 8'h71;    Green = 8'h7d;    Blue = 8'h5a;
end 13'hc13:    begin Red = 8'h6f;    Green = 8'h7a;    Blue = 8'h5e;
end 13'hc14:    begin Red = 8'h72;    Green = 8'h74;    Blue = 8'h55;
end 13'hc15:    begin Red = 8'ha0;    Green = 8'h75;    Blue = 8'h48;
end 13'hc16:    begin Red = 8'h99;    Green = 8'h76;    Blue = 8'h59;
end 13'hc17:    begin Red = 8'h7a;    Green = 8'h72;    Blue = 8'h39;
end 13'hc18:    begin Red = 8'h80;    Green = 8'h78;    Blue = 8'h3f;
end 13'hc19:    begin Red = 8'hce;    Green = 8'hab;    Blue = 8'h84;
end 13'hc1a:    begin Red = 8'hcb;    Green = 8'ha5;    Blue = 8'h87;
end 13'hc1b:    begin Red = 8'hab;    Green = 8'h91;    Blue = 8'h6a;
end 13'hc1c:    begin Red = 8'hd3;    Green = 8'hd7;    Blue = 8'hb7;
end 13'hc1d:    begin Red = 8'ha7;    Green = 8'hae;    Blue = 8'h88;
end 13'hc1e:    begin Red = 8'h85;    Green = 8'h88;    Blue = 8'h71;
end 13'hc1f:    begin Red = 8'hc6;    Green = 8'h8d;    Blue = 8'hba;
end 13'hc20:    begin Red = 8'hbe;    Green = 8'h84;    Blue = 8'hb0;
end 13'hc21:    begin Red = 8'hd5;    Green = 8'he6;    Blue = 8'hdc;
end 13'hc22:    begin Red = 8'hd3;    Green = 8'h9e;    Blue = 8'hc9;
end 13'hc23:    begin Red = 8'hd2;    Green = 8'hdf;    Blue = 8'hde;
end 13'hc24:    begin Red = 8'h9e;    Green = 8'hb1;    Blue = 8'h9c;
end 13'hc25:    begin Red = 8'ha2;    Green = 8'h98;    Blue = 8'h4b;
end 13'hc26:    begin Red = 8'h90;    Green = 8'h8a;    Blue = 8'h4c;
end 13'hc27:    begin Red = 8'h82;    Green = 8'h7b;    Blue = 8'h4f;
end 13'hc28:    begin Red = 8'h81;    Green = 8'h89;    Blue = 8'h45;
end 13'hc29:    begin Red = 8'h80;    Green = 8'h8c;    Blue = 8'h48;
end 13'hc2a:    begin Red = 8'h88;    Green = 8'ha2;    Blue = 8'h48;
end 13'hc2b:    begin Red = 8'h9c;    Green = 8'ha9;    Blue = 8'h85;
end 13'hc2c:    begin Red = 8'h65;    Green = 8'h6c;    Blue = 8'h61;
end 13'hc2d:    begin Red = 8'ha1;    Green = 8'h71;    Blue = 8'h4a;
end 13'hc2e:    begin Red = 8'h7e;    Green = 8'h9f;    Blue = 8'h98;
end 13'hc2f:    begin Red = 8'h7d;    Green = 8'ha1;    Blue = 8'h8a;
end 13'hc30:    begin Red = 8'h7f;    Green = 8'ha2;    Blue = 8'h96;
end 13'hc31:    begin Red = 8'h81;    Green = 8'ha2;    Blue = 8'h9d;
end 13'hc32:    begin Red = 8'h86;    Green = 8'h99;    Blue = 8'h8c;
end 13'hc33:    begin Red = 8'hb1;    Green = 8'h9b;    Blue = 8'h71;
end 13'hc34:    begin Red = 8'hb4;    Green = 8'h97;    Blue = 8'h74;
end 13'hc35:    begin Red = 8'hb7;    Green = 8'h96;    Blue = 8'h76;
end 13'hc36:    begin Red = 8'h9d;    Green = 8'hae;    Blue = 8'h8c;
end 13'hc37:    begin Red = 8'hb3;    Green = 8'hba;    Blue = 8'h94;
end 13'hc38:    begin Red = 8'h9e;    Green = 8'h82;    Blue = 8'h69;
end 13'hc39:    begin Red = 8'hc2;    Green = 8'h7e;    Blue = 8'hb2;
end 13'hc3a:    begin Red = 8'hd6;    Green = 8'h9d;    Blue = 8'hcb;
end 13'hc3b:    begin Red = 8'ha9;    Green = 8'ha3;    Blue = 8'h95;
end 13'hc3c:    begin Red = 8'h93;    Green = 8'h98;    Blue = 8'h4b;
end 13'hc3d:    begin Red = 8'h8f;    Green = 8'h8a;    Blue = 8'h44;
end 13'hc3e:    begin Red = 8'h7f;    Green = 8'h7b;    Blue = 8'h45;
end 13'hc3f:    begin Red = 8'h81;    Green = 8'h7e;    Blue = 8'h4b;
end 13'hc40:    begin Red = 8'h6a;    Green = 8'h6b;    Blue = 8'h50;
end 13'hc41:    begin Red = 8'h86;    Green = 8'ha0;    Blue = 8'h45;
end 13'hc42:    begin Red = 8'h83;    Green = 8'h99;    Blue = 8'h47;
end 13'hc43:    begin Red = 8'h88;    Green = 8'h8f;    Blue = 8'h7e;
end 13'hc44:    begin Red = 8'h7c;    Green = 8'h99;    Blue = 8'h8c;
end 13'hc45:    begin Red = 8'h8c;    Green = 8'h93;    Blue = 8'h85;
end 13'hc46:    begin Red = 8'h7c;    Green = 8'h9c;    Blue = 8'h8e;
end 13'hc47:    begin Red = 8'h98;    Green = 8'h78;    Blue = 8'h49;
end 13'hc48:    begin Red = 8'h77;    Green = 8'h9c;    Blue = 8'h8c;
end 13'hc49:    begin Red = 8'h83;    Green = 8'h9a;    Blue = 8'h82;
end 13'hc4a:    begin Red = 8'hb7;    Green = 8'ha3;    Blue = 8'h78;
end 13'hc4b:    begin Red = 8'hb7;    Green = 8'h94;    Blue = 8'h7f;
end 13'hc4c:    begin Red = 8'ha2;    Green = 8'ha5;    Blue = 8'h8b;
end 13'hc4d:    begin Red = 8'hc1;    Green = 8'h7d;    Blue = 8'haf;
end 13'hc4e:    begin Red = 8'ha3;    Green = 8'hbb;    Blue = 8'haf;
end 13'hc4f:    begin Red = 8'h98;    Green = 8'h8b;    Blue = 8'h42;
end 13'hc50:    begin Red = 8'h93;    Green = 8'h8e;    Blue = 8'h4b;
end 13'hc51:    begin Red = 8'h8d;    Green = 8'h89;    Blue = 8'h48;
end 13'hc52:    begin Red = 8'h75;    Green = 8'h73;    Blue = 8'h4c;
end 13'hc53:    begin Red = 8'h89;    Green = 8'h9d;    Blue = 8'h3e;
end 13'hc54:    begin Red = 8'h81;    Green = 8'h97;    Blue = 8'h3d;
end 13'hc55:    begin Red = 8'h7e;    Green = 8'h90;    Blue = 8'h49;
end 13'hc56:    begin Red = 8'h71;    Green = 8'h77;    Blue = 8'h56;
end 13'hc57:    begin Red = 8'hb5;    Green = 8'h80;    Blue = 8'h5e;
end 13'hc58:    begin Red = 8'h70;    Green = 8'h98;    Blue = 8'h6c;
end 13'hc59:    begin Red = 8'h7d;    Green = 8'haa;    Blue = 8'h78;
end 13'hc5a:    begin Red = 8'h7f;    Green = 8'ha7;    Blue = 8'h76;
end 13'hc5b:    begin Red = 8'h80;    Green = 8'ha5;    Blue = 8'h6c;
end 13'hc5c:    begin Red = 8'hd3;    Green = 8'he0;    Blue = 8'hc1;
end 13'hc5d:    begin Red = 8'he3;    Green = 8'he9;    Blue = 8'hc6;
end 13'hc5e:    begin Red = 8'h6c;    Green = 8'h9a;    Blue = 8'h6b;
end 13'hc5f:    begin Red = 8'h6d;    Green = 8'h93;    Blue = 8'h67;
end 13'hc60:    begin Red = 8'h80;    Green = 8'ha8;    Blue = 8'h70;
end 13'hc61:    begin Red = 8'hbd;    Green = 8'hc2;    Blue = 8'ha3;
end 13'hc62:    begin Red = 8'h90;    Green = 8'ha9;    Blue = 8'he9;
end 13'hc63:    begin Red = 8'hd7;    Green = 8'hdd;    Blue = 8'hbb;
end 13'hc64:    begin Red = 8'hc5;    Green = 8'h82;    Blue = 8'hb1;
end 13'hc65:    begin Red = 8'hc3;    Green = 8'h6c;    Blue = 8'hab;
end 13'hc66:    begin Red = 8'hd6;    Green = 8'he2;    Blue = 8'he0;
end 13'hc67:    begin Red = 8'hcf;    Green = 8'h95;    Blue = 8'hbf;
end 13'hc68:    begin Red = 8'hbd;    Green = 8'hb7;    Blue = 8'ha3;
end 13'hc69:    begin Red = 8'h98;    Green = 8'hb5;    Blue = 8'h8c;
end 13'hc6a:    begin Red = 8'h8b;    Green = 8'h80;    Blue = 8'h34;
end 13'hc6b:    begin Red = 8'h90;    Green = 8'h8c;    Blue = 8'h42;
end 13'hc6c:    begin Red = 8'h88;    Green = 8'h83;    Blue = 8'h45;
end 13'hc6d:    begin Red = 8'h83;    Green = 8'h86;    Blue = 8'h41;
end 13'hc6e:    begin Red = 8'h70;    Green = 8'h71;    Blue = 8'h4a;
end 13'hc6f:    begin Red = 8'h6d;    Green = 8'h6d;    Blue = 8'h52;
end 13'hc70:    begin Red = 8'h88;    Green = 8'ha7;    Blue = 8'h38;
end 13'hc71:    begin Red = 8'h88;    Green = 8'h9d;    Blue = 8'h42;
end 13'hc72:    begin Red = 8'h45;    Green = 8'h3f;    Blue = 8'h3a;
end 13'hc73:    begin Red = 8'h7a;    Green = 8'h91;    Blue = 8'h3d;
end 13'hc74:    begin Red = 8'h46;    Green = 8'h48;    Blue = 8'h3d;
end 13'hc75:    begin Red = 8'h3c;    Green = 8'h3f;    Blue = 8'h37;
end 13'hc76:    begin Red = 8'ha0;    Green = 8'ha6;    Blue = 8'h7d;
end 13'hc77:    begin Red = 8'hae;    Green = 8'h84;    Blue = 8'h5c;
end 13'hc78:    begin Red = 8'h86;    Green = 8'haf;    Blue = 8'h78;
end 13'hc79:    begin Red = 8'h81;    Green = 8'hac;    Blue = 8'h74;
end 13'hc7a:    begin Red = 8'h86;    Green = 8'haa;    Blue = 8'h7d;
end 13'hc7b:    begin Red = 8'hd0;    Green = 8'he1;    Blue = 8'hbe;
end 13'hc7c:    begin Red = 8'he8;    Green = 8'hee;    Blue = 8'hcf;
end 13'hc7d:    begin Red = 8'h73;    Green = 8'h97;    Blue = 8'h69;
end 13'hc7e:    begin Red = 8'h85;    Green = 8'ha7;    Blue = 8'h7b;
end 13'hc7f:    begin Red = 8'h96;    Green = 8'h95;    Blue = 8'h7d;
end 13'hc80:    begin Red = 8'h97;    Green = 8'h9d;    Blue = 8'h80;
end 13'hc81:    begin Red = 8'hc3;    Green = 8'hba;    Blue = 8'hbd;
end 13'hc82:    begin Red = 8'hc0;    Green = 8'hc0;    Blue = 8'hc0;
end 13'hc83:    begin Red = 8'ha0;    Green = 8'h96;    Blue = 8'h48;
end 13'hc84:    begin Red = 8'h9c;    Green = 8'h97;    Blue = 8'h44;
end 13'hc85:    begin Red = 8'h73;    Green = 8'h75;    Blue = 8'h4b;
end 13'hc86:    begin Red = 8'h66;    Green = 8'h68;    Blue = 8'h49;
end 13'hc87:    begin Red = 8'h80;    Green = 8'h94;    Blue = 8'h42;
end 13'hc88:    begin Red = 8'h84;    Green = 8'h9b;    Blue = 8'h43;
end 13'hc89:    begin Red = 8'h85;    Green = 8'h98;    Blue = 8'h42;
end 13'hc8a:    begin Red = 8'h45;    Green = 8'h4c;    Blue = 8'h34;
end 13'hc8b:    begin Red = 8'hb1;    Green = 8'h80;    Blue = 8'h62;
end 13'hc8c:    begin Red = 8'h7e;    Green = 8'h9d;    Blue = 8'h71;
end 13'hc8d:    begin Red = 8'h78;    Green = 8'h96;    Blue = 8'h6d;
end 13'hc8e:    begin Red = 8'h78;    Green = 8'h98;    Blue = 8'h70;
end 13'hc8f:    begin Red = 8'hb7;    Green = 8'hca;    Blue = 8'ha8;
end 13'hc90:    begin Red = 8'hc3;    Green = 8'hc7;    Blue = 8'hab;
end 13'hc91:    begin Red = 8'hd3;    Green = 8'hd9;    Blue = 8'hb4;
end 13'hc92:    begin Red = 8'h98;    Green = 8'h90;    Blue = 8'h68;
end 13'hc93:    begin Red = 8'h7e;    Green = 8'h7d;    Blue = 8'h6c;
end 13'hc94:    begin Red = 8'h9c;    Green = 8'h8d;    Blue = 8'h6d;
end 13'hc95:    begin Red = 8'h90;    Green = 8'h8c;    Blue = 8'h84;
end 13'hc96:    begin Red = 8'ha5;    Green = 8'ha5;    Blue = 8'h88;
end 13'hc97:    begin Red = 8'hf1;    Green = 8'hde;    Blue = 8'hb1;
end 13'hc98:    begin Red = 8'hbf;    Green = 8'h80;    Blue = 8'hb2;
end 13'hc99:    begin Red = 8'hbe;    Green = 8'h75;    Blue = 8'hb3;
end 13'hc9a:    begin Red = 8'hd2;    Green = 8'hd6;    Blue = 8'hd9;
end 13'hc9b:    begin Red = 8'h76;    Green = 8'h69;    Blue = 8'h57;
end 13'hc9c:    begin Red = 8'h78;    Green = 8'h6b;    Blue = 8'h59;
end 13'hc9d:    begin Red = 8'h82;    Green = 8'h75;    Blue = 8'h63;
end 13'hc9e:    begin Red = 8'h83;    Green = 8'h69;    Blue = 8'h5a;
end 13'hc9f:    begin Red = 8'h8b;    Green = 8'h69;    Blue = 8'h5d;
end 13'hca0:    begin Red = 8'ha0;    Green = 8'hbb;    Blue = 8'hb2;
end 13'hca1:    begin Red = 8'h9f;    Green = 8'hc3;    Blue = 8'hc5;
end 13'hca2:    begin Red = 8'h92;    Green = 8'h90;    Blue = 8'h4e;
end 13'hca3:    begin Red = 8'ha6;    Green = 8'ha0;    Blue = 8'h44;
end 13'hca4:    begin Red = 8'ha8;    Green = 8'h9f;    Blue = 8'h46;
end 13'hca5:    begin Red = 8'h8f;    Green = 8'h8f;    Blue = 8'h47;
end 13'hca6:    begin Red = 8'h73;    Green = 8'h71;    Blue = 8'h48;
end 13'hca7:    begin Red = 8'h4f;    Green = 8'h41;    Blue = 8'h4c;
end 13'hca8:    begin Red = 8'h67;    Green = 8'h4a;    Blue = 8'h4c;
end 13'hca9:    begin Red = 8'h78;    Green = 8'h8f;    Blue = 8'h37;
end 13'hcaa:    begin Red = 8'h74;    Green = 8'h75;    Blue = 8'h46;
end 13'hcab:    begin Red = 8'h66;    Green = 8'h55;    Blue = 8'h4c;
end 13'hcac:    begin Red = 8'h42;    Green = 8'h46;    Blue = 8'h35;
end 13'hcad:    begin Red = 8'h82;    Green = 8'h85;    Blue = 8'h68;
end 13'hcae:    begin Red = 8'ha9;    Green = 8'hc4;    Blue = 8'haa;
end 13'hcaf:    begin Red = 8'hb0;    Green = 8'h82;    Blue = 8'h64;
end 13'hcb0:    begin Red = 8'h7f;    Green = 8'ha1;    Blue = 8'h77;
end 13'hcb1:    begin Red = 8'h92;    Green = 8'hbb;    Blue = 8'h86;
end 13'hcb2:    begin Red = 8'h8d;    Green = 8'hb5;    Blue = 8'h84;
end 13'hcb3:    begin Red = 8'he2;    Green = 8'he6;    Blue = 8'hc3;
end 13'hcb4:    begin Red = 8'haa;    Green = 8'haf;    Blue = 8'h90;
end 13'hcb5:    begin Red = 8'ha0;    Green = 8'h7b;    Blue = 8'h5a;
end 13'hcb6:    begin Red = 8'h7b;    Green = 8'h9e;    Blue = 8'h74;
end 13'hcb7:    begin Red = 8'hd5;    Green = 8'hdb;    Blue = 8'hb6;
end 13'hcb8:    begin Red = 8'h9e;    Green = 8'h96;    Blue = 8'h7a;
end 13'hcb9:    begin Red = 8'h92;    Green = 8'h81;    Blue = 8'h7d;
end 13'hcba:    begin Red = 8'hd6;    Green = 8'hda;    Blue = 8'hbe;
end 13'hcbb:    begin Red = 8'hbe;    Green = 8'h7e;    Blue = 8'hb5;
end 13'hcbc:    begin Red = 8'hd5;    Green = 8'hd8;    Blue = 8'hdf;
end 13'hcbd:    begin Red = 8'hd0;    Green = 8'h9b;    Blue = 8'hc6;
end 13'hcbe:    begin Red = 8'h78;    Green = 8'h6f;    Blue = 8'h5d;
end 13'hcbf:    begin Red = 8'h83;    Green = 8'h79;    Blue = 8'h66;
end 13'hcc0:    begin Red = 8'h9b;    Green = 8'hbd;    Blue = 8'hac;
end 13'hcc1:    begin Red = 8'h94;    Green = 8'h87;    Blue = 8'h3b;
end 13'hcc2:    begin Red = 8'h94;    Green = 8'h93;    Blue = 8'h4b;
end 13'hcc3:    begin Red = 8'h53;    Green = 8'h4e;    Blue = 8'h45;
end 13'hcc4:    begin Red = 8'h64;    Green = 8'h57;    Blue = 8'h4d;
end 13'hcc5:    begin Red = 8'h68;    Green = 8'h5d;    Blue = 8'h4e;
end 13'hcc6:    begin Red = 8'h71;    Green = 8'h79;    Blue = 8'h45;
end 13'hcc7:    begin Red = 8'h6b;    Green = 8'h75;    Blue = 8'h43;
end 13'hcc8:    begin Red = 8'h51;    Green = 8'h5b;    Blue = 8'h3b;
end 13'hcc9:    begin Red = 8'h7f;    Green = 8'h8d;    Blue = 8'h65;
end 13'hcca:    begin Red = 8'hac;    Green = 8'h7e;    Blue = 8'h61;
end 13'hccb:    begin Red = 8'hd6;    Green = 8'he4;    Blue = 8'hc6;
end 13'hccc:    begin Red = 8'hde;    Green = 8'he3;    Blue = 8'hc2;
end 13'hccd:    begin Red = 8'h79;    Green = 8'h9c;    Blue = 8'h72;
end 13'hcce:    begin Red = 8'h75;    Green = 8'h83;    Blue = 8'hac;
end 13'hccf:    begin Red = 8'ha7;    Green = 8'h9b;    Blue = 8'h76;
end 13'hcd0:    begin Red = 8'h9c;    Green = 8'h92;    Blue = 8'h71;
end 13'hcd1:    begin Red = 8'hc0;    Green = 8'hc5;    Blue = 8'ha2;
end 13'hcd2:    begin Red = 8'h82;    Green = 8'h78;    Blue = 8'h6b;
end 13'hcd3:    begin Red = 8'h98;    Green = 8'h81;    Blue = 8'h80;
end 13'hcd4:    begin Red = 8'hce;    Green = 8'h98;    Blue = 8'hc5;
end 13'hcd5:    begin Red = 8'hd4;    Green = 8'hd2;    Blue = 8'hdb;
end 13'hcd6:    begin Red = 8'h8c;    Green = 8'h80;    Blue = 8'h6d;
end 13'hcd7:    begin Red = 8'h90;    Green = 8'h83;    Blue = 8'h6e;
end 13'hcd8:    begin Red = 8'h94;    Green = 8'hb2;    Blue = 8'h97;
end 13'hcd9:    begin Red = 8'h7a;    Green = 8'h7a;    Blue = 8'h34;
end 13'hcda:    begin Red = 8'h80;    Green = 8'h85;    Blue = 8'h4a;
end 13'hcdb:    begin Red = 8'h84;    Green = 8'h88;    Blue = 8'h46;
end 13'hcdc:    begin Red = 8'h7d;    Green = 8'h6a;    Blue = 8'h4e;
end 13'hcdd:    begin Red = 8'h67;    Green = 8'h61;    Blue = 8'h4e;
end 13'hcde:    begin Red = 8'h96;    Green = 8'h9d;    Blue = 8'h7b;
end 13'hcdf:    begin Red = 8'hb6;    Green = 8'hc4;    Blue = 8'ha6;
end 13'hce0:    begin Red = 8'h98;    Green = 8'h9c;    Blue = 8'h83;
end 13'hce1:    begin Red = 8'hbb;    Green = 8'hc0;    Blue = 8'h9d;
end 13'hce2:    begin Red = 8'h5c;    Green = 8'h77;    Blue = 8'h9d;
end 13'hce3:    begin Red = 8'h5d;    Green = 8'h78;    Blue = 8'ha0;
end 13'hce4:    begin Red = 8'h5e;    Green = 8'h75;    Blue = 8'ha7;
end 13'hce5:    begin Red = 8'h62;    Green = 8'h74;    Blue = 8'ha3;
end 13'hce6:    begin Red = 8'h8a;    Green = 8'h79;    Blue = 8'h75;
end 13'hce7:    begin Red = 8'h65;    Green = 8'h7e;    Blue = 8'ha7;
end 13'hce8:    begin Red = 8'h6a;    Green = 8'h7e;    Blue = 8'hb3;
end 13'hce9:    begin Red = 8'h65;    Green = 8'h7d;    Blue = 8'hb5;
end 13'hcea:    begin Red = 8'h68;    Green = 8'h85;    Blue = 8'ha8;
end 13'hceb:    begin Red = 8'h8e;    Green = 8'h88;    Blue = 8'h84;
end 13'hcec:    begin Red = 8'h62;    Green = 8'h81;    Blue = 8'haf;
end 13'hced:    begin Red = 8'h8e;    Green = 8'h8f;    Blue = 8'h74;
end 13'hcee:    begin Red = 8'h55;    Green = 8'h78;    Blue = 8'h9e;
end 13'hcef:    begin Red = 8'hd2;    Green = 8'h8d;    Blue = 8'hb7;
end 13'hcf0:    begin Red = 8'hde;    Green = 8'hf1;    Blue = 8'he4;
end 13'hcf1:    begin Red = 8'hd6;    Green = 8'h99;    Blue = 8'hbe;
end 13'hcf2:    begin Red = 8'h87;    Green = 8'h7c;    Blue = 8'h71;
end 13'hcf3:    begin Red = 8'h89;    Green = 8'h7d;    Blue = 8'h6e;
end 13'hcf4:    begin Red = 8'h91;    Green = 8'h79;    Blue = 8'h5d;
end 13'hcf5:    begin Red = 8'ha3;    Green = 8'hb1;    Blue = 8'h9c;
end 13'hcf6:    begin Red = 8'ha4;    Green = 8'hc3;    Blue = 8'hab;
end 13'hcf7:    begin Red = 8'h84;    Green = 8'h7d;    Blue = 8'h34;
end 13'hcf8:    begin Red = 8'h89;    Green = 8'h84;    Blue = 8'h4a;
end 13'hcf9:    begin Red = 8'h8e;    Green = 8'h8c;    Blue = 8'h4d;
end 13'hcfa:    begin Red = 8'h8c;    Green = 8'h74;    Blue = 8'h57;
end 13'hcfb:    begin Red = 8'h78;    Green = 8'h68;    Blue = 8'h4f;
end 13'hcfc:    begin Red = 8'h67;    Green = 8'h5b;    Blue = 8'h4c;
end 13'hcfd:    begin Red = 8'h64;    Green = 8'h5a;    Blue = 8'h4a;
end 13'hcfe:    begin Red = 8'h56;    Green = 8'h61;    Blue = 8'h3f;
end 13'hcff:    begin Red = 8'h8b;    Green = 8'h90;    Blue = 8'h6f;
end 13'hd00:    begin Red = 8'h68;    Green = 8'h6d;    Blue = 8'h44;
end 13'hd01:    begin Red = 8'haa;    Green = 8'hc2;    Blue = 8'ha7;
end 13'hd02:    begin Red = 8'hab;    Green = 8'hbe;    Blue = 8'h9f;
end 13'hd03:    begin Red = 8'haa;    Green = 8'h80;    Blue = 8'h59;
end 13'hd04:    begin Red = 8'h8d;    Green = 8'hc2;    Blue = 8'h89;
end 13'hd05:    begin Red = 8'h8e;    Green = 8'hbb;    Blue = 8'h85;
end 13'hd06:    begin Red = 8'h8b;    Green = 8'hbb;    Blue = 8'h88;
end 13'hd07:    begin Red = 8'h95;    Green = 8'h9a;    Blue = 8'h7f;
end 13'hd08:    begin Red = 8'ha3;    Green = 8'h7d;    Blue = 8'h5c;
end 13'hd09:    begin Red = 8'ha5;    Green = 8'h86;    Blue = 8'h64;
end 13'hd0a:    begin Red = 8'h76;    Green = 8'h9f;    Blue = 8'h71;
end 13'hd0b:    begin Red = 8'h97;    Green = 8'h8d;    Blue = 8'h7a;
end 13'hd0c:    begin Red = 8'h80;    Green = 8'h7e;    Blue = 8'h72;
end 13'hd0d:    begin Red = 8'ha5;    Green = 8'h90;    Blue = 8'h87;
end 13'hd0e:    begin Red = 8'hd0;    Green = 8'hd9;    Blue = 8'hbb;
end 13'hd0f:    begin Red = 8'h97;    Green = 8'h85;    Blue = 8'h7b;
end 13'hd10:    begin Red = 8'hbb;    Green = 8'h75;    Blue = 8'ha4;
end 13'hd11:    begin Red = 8'hce;    Green = 8'hdb;    Blue = 8'hdb;
end 13'hd12:    begin Red = 8'hcd;    Green = 8'h8c;    Blue = 8'hc0;
end 13'hd13:    begin Red = 8'hc8;    Green = 8'h9d;    Blue = 8'hc4;
end 13'hd14:    begin Red = 8'ha0;    Green = 8'h92;    Blue = 8'h7d;
end 13'hd15:    begin Red = 8'hb5;    Green = 8'hb0;    Blue = 8'ha3;
end 13'hd16:    begin Red = 8'ha1;    Green = 8'hbb;    Blue = 8'ha8;
end 13'hd17:    begin Red = 8'h73;    Green = 8'h7e;    Blue = 8'h3f;
end 13'hd18:    begin Red = 8'h57;    Green = 8'h4b;    Blue = 8'h3a;
end 13'hd19:    begin Red = 8'h7c;    Green = 8'h66;    Blue = 8'h4f;
end 13'hd1a:    begin Red = 8'h7a;    Green = 8'h6c;    Blue = 8'h4f;
end 13'hd1b:    begin Red = 8'h75;    Green = 8'h65;    Blue = 8'h51;
end 13'hd1c:    begin Red = 8'h4b;    Green = 8'h46;    Blue = 8'h3b;
end 13'hd1d:    begin Red = 8'h50;    Green = 8'h4b;    Blue = 8'h38;
end 13'hd1e:    begin Red = 8'h71;    Green = 8'h7b;    Blue = 8'h65;
end 13'hd1f:    begin Red = 8'haf;    Green = 8'h96;    Blue = 8'h7f;
end 13'hd20:    begin Red = 8'h75;    Green = 8'h78;    Blue = 8'h66;
end 13'hd21:    begin Red = 8'h9d;    Green = 8'ha2;    Blue = 8'h84;
end 13'hd22:    begin Red = 8'hcb;    Green = 8'hb5;    Blue = 8'h90;
end 13'hd23:    begin Red = 8'hce;    Green = 8'hb9;    Blue = 8'h97;
end 13'hd24:    begin Red = 8'hb7;    Green = 8'h75;    Blue = 8'ha8;
end 13'hd25:    begin Red = 8'hcb;    Green = 8'h96;    Blue = 8'hc1;
end 13'hd26:    begin Red = 8'h96;    Green = 8'h88;    Blue = 8'h78;
end 13'hd27:    begin Red = 8'hde;    Green = 8'hd8;    Blue = 8'hc7;
end 13'hd28:    begin Red = 8'h94;    Green = 8'h86;    Blue = 8'h76;
end 13'hd29:    begin Red = 8'he6;    Green = 8'he3;    Blue = 8'hcf;
end 13'hd2a:    begin Red = 8'ha3;    Green = 8'hb8;    Blue = 8'h94;
end 13'hd2b:    begin Red = 8'h55;    Green = 8'h4e;    Blue = 8'h42;
end 13'hd2c:    begin Red = 8'h5a;    Green = 8'h51;    Blue = 8'h41;
end 13'hd2d:    begin Red = 8'h6f;    Green = 8'h63;    Blue = 8'h49;
end 13'hd2e:    begin Red = 8'h71;    Green = 8'h63;    Blue = 8'h4d;
end 13'hd2f:    begin Red = 8'h75;    Green = 8'h6a;    Blue = 8'h4d;
end 13'hd30:    begin Red = 8'h72;    Green = 8'h61;    Blue = 8'h49;
end 13'hd31:    begin Red = 8'h56;    Green = 8'h52;    Blue = 8'h3b;
end 13'hd32:    begin Red = 8'h69;    Green = 8'h66;    Blue = 8'h46;
end 13'hd33:    begin Red = 8'h61;    Green = 8'h57;    Blue = 8'h37;
end 13'hd34:    begin Red = 8'hcd;    Green = 8'hdb;    Blue = 8'hbb;
end 13'hd35:    begin Red = 8'ha8;    Green = 8'hac;    Blue = 8'h90;
end 13'hd36:    begin Red = 8'hcf;    Green = 8'hbb;    Blue = 8'h9b;
end 13'hd37:    begin Red = 8'ha7;    Green = 8'hc2;    Blue = 8'ha9;
end 13'hd38:    begin Red = 8'h7f;    Green = 8'h70;    Blue = 8'h55;
end 13'hd39:    begin Red = 8'h6e;    Green = 8'h61;    Blue = 8'h47;
end 13'hd3a:    begin Red = 8'h60;    Green = 8'h5d;    Blue = 8'h42;
end 13'hd3b:    begin Red = 8'ha9;    Green = 8'hc9;    Blue = 8'had;
end 13'hd3c:    begin Red = 8'ha8;    Green = 8'hb2;    Blue = 8'h92;
end 13'hd3d:    begin Red = 8'h71;    Green = 8'h90;    Blue = 8'h7c;
end 13'hd3e:    begin Red = 8'hd8;    Green = 8'he6;    Blue = 8'hc7;
end 13'hd3f:    begin Red = 8'hbf;    Green = 8'ha8;    Blue = 8'h88;
end 13'hd40:    begin Red = 8'hb9;    Green = 8'ha8;    Blue = 8'h86;
end 13'hd41:    begin Red = 8'hc2;    Green = 8'ha8;    Blue = 8'h8a;
end 13'hd42:    begin Red = 8'hc3;    Green = 8'hb9;    Blue = 8'hc7;
end 13'hd43:    begin Red = 8'hbb;    Green = 8'h86;    Blue = 8'haf;
end 13'hd44:    begin Red = 8'haf;    Green = 8'h74;    Blue = 8'ha3;
end 13'hd45:    begin Red = 8'hd6;    Green = 8'he0;    Blue = 8'hd2;
end 13'hd46:    begin Red = 8'hce;    Green = 8'h93;    Blue = 8'hba;
end 13'hd47:    begin Red = 8'h79;    Green = 8'h5e;    Blue = 8'h42;
end 13'hd48:    begin Red = 8'h74;    Green = 8'h62;    Blue = 8'h43;
end 13'hd49:    begin Red = 8'h92;    Green = 8'h72;    Blue = 8'h55;
end 13'hd4a:    begin Red = 8'h83;    Green = 8'h6a;    Blue = 8'h51;
end 13'hd4b:    begin Red = 8'h8d;    Green = 8'h72;    Blue = 8'h55;
end 13'hd4c:    begin Red = 8'h48;    Green = 8'h4a;    Blue = 8'h3b;
end 13'hd4d:    begin Red = 8'h53;    Green = 8'h50;    Blue = 8'h34;
end 13'hd4e:    begin Red = 8'hb7;    Green = 8'hc0;    Blue = 8'h9a;
end 13'hd4f:    begin Red = 8'h47;    Green = 8'h3f;    Blue = 8'h40;
end 13'hd50:    begin Red = 8'h52;    Green = 8'h4a;    Blue = 8'h45;
end 13'hd51:    begin Red = 8'h8c;    Green = 8'h86;    Blue = 8'h70;
end 13'hd52:    begin Red = 8'hc3;    Green = 8'hc9;    Blue = 8'ha6;
end 13'hd53:    begin Red = 8'h4e;    Green = 8'h44;    Blue = 8'h47;
end 13'hd54:    begin Red = 8'he9;    Green = 8'hd0;    Blue = 8'hab;
end 13'hd55:    begin Red = 8'hbb;    Green = 8'hc4;    Blue = 8'hc1;
end 13'hd56:    begin Red = 8'hce;    Green = 8'hd3;    Blue = 8'hd0;
end 13'hd57:    begin Red = 8'h96;    Green = 8'h84;    Blue = 8'h77;
end 13'hd58:    begin Red = 8'he8;    Green = 8'he5;    Blue = 8'hd1;
end 13'hd59:    begin Red = 8'hea;    Green = 8'hae;    Blue = 8'h80;
end 13'hd5a:    begin Red = 8'he6;    Green = 8'hae;    Blue = 8'h84;
end 13'hd5b:    begin Red = 8'he9;    Green = 8'haf;    Blue = 8'h86;
end 13'hd5c:    begin Red = 8'he5;    Green = 8'had;    Blue = 8'h7c;
end 13'hd5d:    begin Red = 8'hfc;    Green = 8'hb6;    Blue = 8'h96;
end 13'hd5e:    begin Red = 8'hff;    Green = 8'hb7;    Blue = 8'h92;
end 13'hd5f:    begin Red = 8'h5d;    Green = 8'h77;    Blue = 8'h38;
end 13'hd60:    begin Red = 8'h8c;    Green = 8'h73;    Blue = 8'h52;
end 13'hd61:    begin Red = 8'h7f;    Green = 8'h69;    Blue = 8'h4a;
end 13'hd62:    begin Red = 8'h68;    Green = 8'h5d;    Blue = 8'h3f;
end 13'hd63:    begin Red = 8'h84;    Green = 8'h69;    Blue = 8'h4a;
end 13'hd64:    begin Red = 8'haf;    Green = 8'hc2;    Blue = 8'h9a;
end 13'hd65:    begin Red = 8'h74;    Green = 8'h61;    Blue = 8'h59;
end 13'hd66:    begin Red = 8'h77;    Green = 8'h61;    Blue = 8'h5c;
end 13'hd67:    begin Red = 8'hcf;    Green = 8'hde;    Blue = 8'hbc;
end 13'hd68:    begin Red = 8'hda;    Green = 8'hdf;    Blue = 8'hbb;
end 13'hd69:    begin Red = 8'hbb;    Green = 8'hb3;    Blue = 8'hc1;
end 13'hd6a:    begin Red = 8'h86;    Green = 8'haa;    Blue = 8'h8b;
end 13'hd6b:    begin Red = 8'hf3;    Green = 8'hac;    Blue = 8'h89;
end 13'hd6c:    begin Red = 8'hff;    Green = 8'hb3;    Blue = 8'h8e;
end 13'hd6d:    begin Red = 8'hf9;    Green = 8'hbb;    Blue = 8'h8d;
end 13'hd6e:    begin Red = 8'h5a;    Green = 8'h76;    Blue = 8'h3d;
end 13'hd6f:    begin Red = 8'he3;    Green = 8'hb1;    Blue = 8'h87;
end 13'hd70:    begin Red = 8'h90;    Green = 8'h6e;    Blue = 8'h4d;
end 13'hd71:    begin Red = 8'h70;    Green = 8'h64;    Blue = 8'h45;
end 13'hd72:    begin Red = 8'h72;    Green = 8'h65;    Blue = 8'h42;
end 13'hd73:    begin Red = 8'h7c;    Green = 8'h6b;    Blue = 8'h47;
end 13'hd74:    begin Red = 8'h6c;    Green = 8'h65;    Blue = 8'h42;
end 13'hd75:    begin Red = 8'h6f;    Green = 8'h63;    Blue = 8'h42;
end 13'hd76:    begin Red = 8'h88;    Green = 8'h69;    Blue = 8'h4c;
end 13'hd77:    begin Red = 8'h84;    Green = 8'h90;    Blue = 8'h74;
end 13'hd78:    begin Red = 8'h78;    Green = 8'h63;    Blue = 8'h55;
end 13'hd79:    begin Red = 8'h75;    Green = 8'h68;    Blue = 8'h54;
end 13'hd7a:    begin Red = 8'hdb;    Green = 8'he2;    Blue = 8'hbc;
end 13'hd7b:    begin Red = 8'h7c;    Green = 8'h71;    Blue = 8'h62;
end 13'hd7c:    begin Red = 8'hbe;    Green = 8'hc4;    Blue = 8'ha7;
end 13'hd7d:    begin Red = 8'h9d;    Green = 8'h9f;    Blue = 8'h81;
end 13'hd7e:    begin Red = 8'he9;    Green = 8'hd2;    Blue = 8'hb3;
end 13'hd7f:    begin Red = 8'hb7;    Green = 8'h83;    Blue = 8'hae;
end 13'hd80:    begin Red = 8'hb5;    Green = 8'h79;    Blue = 8'ha6;
end 13'hd81:    begin Red = 8'hcc;    Green = 8'h8c;    Blue = 8'hb8;
end 13'hd82:    begin Red = 8'hbe;    Green = 8'h88;    Blue = 8'had;
end 13'hd83:    begin Red = 8'hd6;    Green = 8'hdd;    Blue = 8'hc7;
end 13'hd84:    begin Red = 8'h9f;    Green = 8'hb3;    Blue = 8'h90;
end 13'hd85:    begin Red = 8'hff;    Green = 8'haa;    Blue = 8'h80;
end 13'hd86:    begin Red = 8'he6;    Green = 8'hac;    Blue = 8'h88;
end 13'hd87:    begin Red = 8'hd2;    Green = 8'h9c;    Blue = 8'h73;
end 13'hd88:    begin Red = 8'heb;    Green = 8'hb1;    Blue = 8'h87;
end 13'hd89:    begin Red = 8'hd6;    Green = 8'ha0;    Blue = 8'h77;
end 13'hd8a:    begin Red = 8'hea;    Green = 8'had;    Blue = 8'h84;
end 13'hd8b:    begin Red = 8'hed;    Green = 8'hb0;    Blue = 8'h82;
end 13'hd8c:    begin Red = 8'heb;    Green = 8'ha9;    Blue = 8'h7e;
end 13'hd8d:    begin Red = 8'hea;    Green = 8'hb3;    Blue = 8'h84;
end 13'hd8e:    begin Red = 8'h63;    Green = 8'h54;    Blue = 8'h3a;
end 13'hd8f:    begin Red = 8'h78;    Green = 8'h66;    Blue = 8'h49;
end 13'hd90:    begin Red = 8'h4d;    Green = 8'h5b;    Blue = 8'h50;
end 13'hd91:    begin Red = 8'hbd;    Green = 8'h88;    Blue = 8'h62;
end 13'hd92:    begin Red = 8'h75;    Green = 8'h69;    Blue = 8'h46;
end 13'hd93:    begin Red = 8'h77;    Green = 8'h65;    Blue = 8'h44;
end 13'hd94:    begin Red = 8'h71;    Green = 8'h60;    Blue = 8'h41;
end 13'hd95:    begin Red = 8'he7;    Green = 8'hf6;    Blue = 8'hcf;
end 13'hd96:    begin Red = 8'hce;    Green = 8'hdb;    Blue = 8'hb0;
end 13'hd97:    begin Red = 8'hd4;    Green = 8'he2;    Blue = 8'hc4;
end 13'hd98:    begin Red = 8'hd5;    Green = 8'hd9;    Blue = 8'hbb;
end 13'hd99:    begin Red = 8'hb4;    Green = 8'h80;    Blue = 8'had;
end 13'hd9a:    begin Red = 8'hb6;    Green = 8'h6e;    Blue = 8'h98;
end 13'hd9b:    begin Red = 8'hd8;    Green = 8'he1;    Blue = 8'hde;
end 13'hd9c:    begin Red = 8'hde;    Green = 8'he6;    Blue = 8'hde;
end 13'hd9d:    begin Red = 8'hda;    Green = 8'hea;    Blue = 8'he1;
end 13'hd9e:    begin Red = 8'hd3;    Green = 8'h93;    Blue = 8'h61;
end 13'hd9f:    begin Red = 8'hd2;    Green = 8'h8f;    Blue = 8'h5f;
end 13'hda0:    begin Red = 8'hfd;    Green = 8'hb3;    Blue = 8'h85;
end 13'hda1:    begin Red = 8'hff;    Green = 8'hb8;    Blue = 8'h88;
end 13'hda2:    begin Red = 8'hed;    Green = 8'ha5;    Blue = 8'h74;
end 13'hda3:    begin Red = 8'hf9;    Green = 8'hb2;    Blue = 8'h7d;
end 13'hda4:    begin Red = 8'hf9;    Green = 8'hb2;    Blue = 8'h82;
end 13'hda5:    begin Red = 8'hfb;    Green = 8'hb7;    Blue = 8'h86;
end 13'hda6:    begin Red = 8'hf3;    Green = 8'hb0;    Blue = 8'h7d;
end 13'hda7:    begin Red = 8'hf9;    Green = 8'hac;    Blue = 8'h7e;
end 13'hda8:    begin Red = 8'hf5;    Green = 8'hab;    Blue = 8'h7c;
end 13'hda9:    begin Red = 8'he8;    Green = 8'ha2;    Blue = 8'h6f;
end 13'hdaa:    begin Red = 8'he7;    Green = 8'ha4;    Blue = 8'h71;
end 13'hdab:    begin Red = 8'hde;    Green = 8'h9b;    Blue = 8'h6b;
end 13'hdac:    begin Red = 8'hfc;    Green = 8'haf;    Blue = 8'h81;
end 13'hdad:    begin Red = 8'hfd;    Green = 8'ha9;    Blue = 8'h83;
end 13'hdae:    begin Red = 8'hfe;    Green = 8'hac;    Blue = 8'h71;
end 13'hdaf:    begin Red = 8'hfb;    Green = 8'hab;    Blue = 8'h75;
end 13'hdb0:    begin Red = 8'he7;    Green = 8'had;    Blue = 8'h81;
end 13'hdb1:    begin Red = 8'hd2;    Green = 8'h99;    Blue = 8'h70;
end 13'hdb2:    begin Red = 8'hce;    Green = 8'h96;    Blue = 8'h6c;
end 13'hdb3:    begin Red = 8'hee;    Green = 8'hb4;    Blue = 8'h8a;
end 13'hdb4:    begin Red = 8'hf0;    Green = 8'hac;    Blue = 8'h80;
end 13'hdb5:    begin Red = 8'hf7;    Green = 8'hb6;    Blue = 8'h89;
end 13'hdb6:    begin Red = 8'hfa;    Green = 8'hc0;    Blue = 8'h98;
end 13'hdb7:    begin Red = 8'h74;    Green = 8'h69;    Blue = 8'h51;
end 13'hdb8:    begin Red = 8'h74;    Green = 8'h68;    Blue = 8'h49;
end 13'hdb9:    begin Red = 8'h4e;    Green = 8'h5a;    Blue = 8'h4c;
end 13'hdba:    begin Red = 8'hc7;    Green = 8'h8f;    Blue = 8'h65;
end 13'hdbb:    begin Red = 8'hd6;    Green = 8'h90;    Blue = 8'h6b;
end 13'hdbc:    begin Red = 8'hde;    Green = 8'h96;    Blue = 8'h6c;
end 13'hdbd:    begin Red = 8'h71;    Green = 8'h6e;    Blue = 8'h55;
end 13'hdbe:    begin Red = 8'h5c;    Green = 8'h59;    Blue = 8'h34;
end 13'hdbf:    begin Red = 8'hd4;    Green = 8'h94;    Blue = 8'h64;
end 13'hdc0:    begin Red = 8'hbe;    Green = 8'hd2;    Blue = 8'hac;
end 13'hdc1:    begin Red = 8'hbe;    Green = 8'hbc;    Blue = 8'h9b;
end 13'hdc2:    begin Red = 8'hbb;    Green = 8'hca;    Blue = 8'hac;
end 13'hdc3:    begin Red = 8'he3;    Green = 8'hc7;    Blue = 8'ha9;
end 13'hdc4:    begin Red = 8'hb7;    Green = 8'ha8;    Blue = 8'h8c;
end 13'hdc5:    begin Red = 8'he2;    Green = 8'hce;    Blue = 8'hb5;
end 13'hdc6:    begin Red = 8'he7;    Green = 8'hcb;    Blue = 8'hb2;
end 13'hdc7:    begin Red = 8'hb2;    Green = 8'h82;    Blue = 8'hac;
end 13'hdc8:    begin Red = 8'hb2;    Green = 8'h6f;    Blue = 8'ha0;
end 13'hdc9:    begin Red = 8'he9;    Green = 8'hb3;    Blue = 8'h7a;
end 13'hdca:    begin Red = 8'h90;    Green = 8'hb4;    Blue = 8'h9d;
end 13'hdcb:    begin Red = 8'hf0;    Green = 8'haa;    Blue = 8'h84;
end 13'hdcc:    begin Red = 8'h64;    Green = 8'h62;    Blue = 8'h50;
end 13'hdcd:    begin Red = 8'h4d;    Green = 8'h59;    Blue = 8'h48;
end 13'hdce:    begin Red = 8'h76;    Green = 8'h6c;    Blue = 8'h52;
end 13'hdcf:    begin Red = 8'hc0;    Green = 8'hd2;    Blue = 8'hb5;
end 13'hdd0:    begin Red = 8'h98;    Green = 8'h94;    Blue = 8'h75;
end 13'hdd1:    begin Red = 8'hc7;    Green = 8'hcc;    Blue = 8'hae;
end 13'hdd2:    begin Red = 8'hfd;    Green = 8'he5;    Blue = 8'hb9;
end 13'hdd3:    begin Red = 8'h6b;    Green = 8'h5a;    Blue = 8'h56;
end 13'hdd4:    begin Red = 8'hf6;    Green = 8'he6;    Blue = 8'hb4;
end 13'hdd5:    begin Red = 8'hff;    Green = 8'he7;    Blue = 8'hb4;
end 13'hdd6:    begin Red = 8'hf9;    Green = 8'he5;    Blue = 8'hb6;
end 13'hdd7:    begin Red = 8'haf;    Green = 8'h80;    Blue = 8'ha8;
end 13'hdd8:    begin Red = 8'hae;    Green = 8'h6b;    Blue = 8'h9c;
end 13'hdd9:    begin Red = 8'hc0;    Green = 8'h8d;    Blue = 8'hb7;
end 13'hdda:    begin Red = 8'hd1;    Green = 8'h98;    Blue = 8'h6d;
end 13'hddb:    begin Red = 8'he3;    Green = 8'hae;    Blue = 8'h8a;
end 13'hddc:    begin Red = 8'he7;    Green = 8'haf;    Blue = 8'h7d;
end 13'hddd:    begin Red = 8'hee;    Green = 8'hab;    Blue = 8'h8d;
end 13'hdde:    begin Red = 8'h84;    Green = 8'hba;    Blue = 8'h9e;
end 13'hddf:    begin Red = 8'hd0;    Green = 8'ha6;    Blue = 8'h7b;
end 13'hde0:    begin Red = 8'hd6;    Green = 8'ha7;    Blue = 8'h7c;
end 13'hde1:    begin Red = 8'h80;    Green = 8'h88;    Blue = 8'h67;
end 13'hde2:    begin Red = 8'h86;    Green = 8'h90;    Blue = 8'h69;
end 13'hde3:    begin Red = 8'hc7;    Green = 8'h8c;    Blue = 8'h67;
end 13'hde4:    begin Red = 8'hc3;    Green = 8'h8d;    Blue = 8'h64;
end 13'hde5:    begin Red = 8'hc4;    Green = 8'h89;    Blue = 8'h62;
end 13'hde6:    begin Red = 8'hd8;    Green = 8'he8;    Blue = 8'hcc;
end 13'hde7:    begin Red = 8'ha6;    Green = 8'hae;    Blue = 8'h92;
end 13'hde8:    begin Red = 8'h9b;    Green = 8'had;    Blue = 8'h9c;
end 13'hde9:    begin Red = 8'hca;    Green = 8'h88;    Blue = 8'h65;
end 13'hdea:    begin Red = 8'h5e;    Green = 8'h52;    Blue = 8'h50;
end 13'hdeb:    begin Red = 8'h61;    Green = 8'h52;    Blue = 8'h4e;
end 13'hdec:    begin Red = 8'h5e;    Green = 8'h53;    Blue = 8'h4a;
end 13'hded:    begin Red = 8'ha5;    Green = 8'ha9;    Blue = 8'h89;
end 13'hdee:    begin Red = 8'h5c;    Green = 8'h55;    Blue = 8'h4e;
end 13'hdef:    begin Red = 8'hf5;    Green = 8'he0;    Blue = 8'hb1;
end 13'hdf0:    begin Red = 8'hcf;    Green = 8'h9a;    Blue = 8'h71;
end 13'hdf1:    begin Red = 8'he1;    Green = 8'hb4;    Blue = 8'h84;
end 13'hdf2:    begin Red = 8'he7;    Green = 8'hb4;    Blue = 8'h83;
end 13'hdf3:    begin Red = 8'h7d;    Green = 8'hba;    Blue = 8'h9f;
end 13'hdf4:    begin Red = 8'h8e;    Green = 8'hb5;    Blue = 8'ha3;
end 13'hdf5:    begin Red = 8'hf1;    Green = 8'ha8;    Blue = 8'h89;
end 13'hdf6:    begin Red = 8'hd6;    Green = 8'hac;    Blue = 8'h80;
end 13'hdf7:    begin Red = 8'he1;    Green = 8'hac;    Blue = 8'h82;
end 13'hdf8:    begin Red = 8'h86;    Green = 8'h8b;    Blue = 8'h68;
end 13'hdf9:    begin Red = 8'h5e;    Green = 8'h68;    Blue = 8'h56;
end 13'hdfa:    begin Red = 8'h3f;    Green = 8'h52;    Blue = 8'h43;
end 13'hdfb:    begin Red = 8'hc4;    Green = 8'h90;    Blue = 8'h61;
end 13'hdfc:    begin Red = 8'hcb;    Green = 8'h8d;    Blue = 8'h5c;
end 13'hdfd:    begin Red = 8'hbf;    Green = 8'h8d;    Blue = 8'h65;
end 13'hdfe:    begin Red = 8'hdc;    Green = 8'hec;    Blue = 8'hd0;
end 13'hdff:    begin Red = 8'h94;    Green = 8'hbe;    Blue = 8'ha6;
end 13'he00:    begin Red = 8'ha1;    Green = 8'haf;    Blue = 8'h8b;
end 13'he01:    begin Red = 8'h93;    Green = 8'h8c;    Blue = 8'h82;
end 13'he02:    begin Red = 8'ha3;    Green = 8'h6c;    Blue = 8'h97;
end 13'he03:    begin Red = 8'hc0;    Green = 8'h8a;    Blue = 8'haf;
end 13'he04:    begin Red = 8'hd4;    Green = 8'h9f;    Blue = 8'h75;
end 13'he05:    begin Red = 8'ha4;    Green = 8'hb2;    Blue = 8'h98;
end 13'he06:    begin Red = 8'he4;    Green = 8'haa;    Blue = 8'h80;
end 13'he07:    begin Red = 8'hbb;    Green = 8'h8c;    Blue = 8'h65;
end 13'he08:    begin Red = 8'hbc;    Green = 8'hce;    Blue = 8'haf;
end 13'he09:    begin Red = 8'hd2;    Green = 8'h81;    Blue = 8'h4a;
end 13'he0a:    begin Red = 8'h88;    Green = 8'hd9;    Blue = 8'hf4;
end 13'he0b:    begin Red = 8'hb9;    Green = 8'hbe;    Blue = 8'h9b;
end 13'he0c:    begin Red = 8'h5e;    Green = 8'h77;    Blue = 8'ha3;
end 13'he0d:    begin Red = 8'h5b;    Green = 8'h76;    Blue = 8'ha9;
end 13'he0e:    begin Red = 8'h94;    Green = 8'ha9;    Blue = 8'hfd;
end 13'he0f:    begin Red = 8'hf8;    Green = 8'he0;    Blue = 8'hb5;
end 13'he10:    begin Red = 8'h5e;    Green = 8'h73;    Blue = 8'hae;
end 13'he11:    begin Red = 8'h96;    Green = 8'hb1;    Blue = 8'hff;
end 13'he12:    begin Red = 8'h95;    Green = 8'h7f;    Blue = 8'h75;
end 13'he13:    begin Red = 8'ha7;    Green = 8'h78;    Blue = 8'ha1;
end 13'he14:    begin Red = 8'hbb;    Green = 8'h80;    Blue = 8'had;
end 13'he15:    begin Red = 8'hb5;    Green = 8'h7c;    Blue = 8'hae;
end 13'he16:    begin Red = 8'hbe;    Green = 8'h6c;    Blue = 8'ha7;
end 13'he17:    begin Red = 8'h88;    Green = 8'hc0;    Blue = 8'ha5;
end 13'he18:    begin Red = 8'hca;    Green = 8'h92;    Blue = 8'h69;
end 13'he19:    begin Red = 8'he5;    Green = 8'ha9;    Blue = 8'h7d;
end 13'he1a:    begin Red = 8'hc0;    Green = 8'h82;    Blue = 8'h5b;
end 13'he1b:    begin Red = 8'hb8;    Green = 8'h8a;    Blue = 8'h64;
end 13'he1c:    begin Red = 8'hca;    Green = 8'h8d;    Blue = 8'h65;
end 13'he1d:    begin Red = 8'hca;    Green = 8'h87;    Blue = 8'h5b;
end 13'he1e:    begin Red = 8'hd3;    Green = 8'h80;    Blue = 8'h4e;
end 13'he1f:    begin Red = 8'h8a;    Green = 8'hd6;    Blue = 8'hf8;
end 13'he20:    begin Red = 8'h67;    Green = 8'h73;    Blue = 8'ha2;
end 13'he21:    begin Red = 8'h65;    Green = 8'h75;    Blue = 8'ha7;
end 13'he22:    begin Red = 8'h8c;    Green = 8'hb7;    Blue = 8'hff;
end 13'he23:    begin Red = 8'he1;    Green = 8'hce;    Blue = 8'ha9;
end 13'he24:    begin Red = 8'h5e;    Green = 8'h71;    Blue = 8'ha9;
end 13'he25:    begin Red = 8'h60;    Green = 8'h7b;    Blue = 8'hac;
end 13'he26:    begin Red = 8'h85;    Green = 8'hb2;    Blue = 8'hf4;
end 13'he27:    begin Red = 8'hac;    Green = 8'h6e;    Blue = 8'ha4;
end 13'he28:    begin Red = 8'ha7;    Green = 8'h68;    Blue = 8'h98;
end 13'he29:    begin Red = 8'hbb;    Green = 8'h7a;    Blue = 8'hac;
end 13'he2a:    begin Red = 8'hb2;    Green = 8'h73;    Blue = 8'ha7;
end 13'he2b:    begin Red = 8'hc5;    Green = 8'h8c;    Blue = 8'h61;
end 13'he2c:    begin Red = 8'hf2;    Green = 8'hb6;    Blue = 8'h8c;
end 13'he2d:    begin Red = 8'h7d;    Green = 8'hbb;    Blue = 8'ha7;
end 13'he2e:    begin Red = 8'h94;    Green = 8'hb5;    Blue = 8'h9d;
end 13'he2f:    begin Red = 8'h88;    Green = 8'hb6;    Blue = 8'h9c;
end 13'he30:    begin Red = 8'he8;    Green = 8'hb2;    Blue = 8'h81;
end 13'he31:    begin Red = 8'hc1;    Green = 8'h8c;    Blue = 8'h62;
end 13'he32:    begin Red = 8'hc6;    Green = 8'h92;    Blue = 8'h67;
end 13'he33:    begin Red = 8'hbe;    Green = 8'h87;    Blue = 8'h5d;
end 13'he34:    begin Red = 8'hc3;    Green = 8'h87;    Blue = 8'h5f;
end 13'he35:    begin Red = 8'hd6;    Green = 8'hea;    Blue = 8'hcd;
end 13'he36:    begin Red = 8'hc5;    Green = 8'h85;    Blue = 8'h5d;
end 13'he37:    begin Red = 8'hc7;    Green = 8'h89;    Blue = 8'h60;
end 13'he38:    begin Red = 8'hc6;    Green = 8'h87;    Blue = 8'h5a;
end 13'he39:    begin Red = 8'hbb;    Green = 8'h8b;    Blue = 8'h60;
end 13'he3a:    begin Red = 8'h74;    Green = 8'he7;    Blue = 8'hff;
end 13'he3b:    begin Red = 8'h7d;    Green = 8'hd9;    Blue = 8'hf8;
end 13'he3c:    begin Red = 8'h7b;    Green = 8'hd5;    Blue = 8'hf5;
end 13'he3d:    begin Red = 8'h79;    Green = 8'hd6;    Blue = 8'hf2;
end 13'he3e:    begin Red = 8'h81;    Green = 8'hd6;    Blue = 8'hf8;
end 13'he3f:    begin Red = 8'h80;    Green = 8'he1;    Blue = 8'hff;
end 13'he40:    begin Red = 8'hb6;    Green = 8'h9b;    Blue = 8'h7b;
end 13'he41:    begin Red = 8'hd4;    Green = 8'hde;    Blue = 8'hbc;
end 13'he42:    begin Red = 8'h8c;    Green = 8'h77;    Blue = 8'h69;
end 13'he43:    begin Red = 8'h98;    Green = 8'h85;    Blue = 8'h7f;
end 13'he44:    begin Red = 8'heb;    Green = 8'ha8;    Blue = 8'h85;
end 13'he45:    begin Red = 8'hf0;    Green = 8'hab;    Blue = 8'h88;
end 13'he46:    begin Red = 8'he3;    Green = 8'haf;    Blue = 8'h7f;
end 13'he47:    begin Red = 8'h92;    Green = 8'hb3;    Blue = 8'ha3;
end 13'he48:    begin Red = 8'he4;    Green = 8'hac;    Blue = 8'h75;
end 13'he49:    begin Red = 8'hc9;    Green = 8'h90;    Blue = 8'h67;
end 13'he4a:    begin Red = 8'hd0;    Green = 8'he2;    Blue = 8'hc5;
end 13'he4b:    begin Red = 8'hd9;    Green = 8'h9c;    Blue = 8'h73;
end 13'he4c:    begin Red = 8'hcc;    Green = 8'h97;    Blue = 8'h75;
end 13'he4d:    begin Red = 8'hca;    Green = 8'h93;    Blue = 8'h74;
end 13'he4e:    begin Red = 8'hca;    Green = 8'h95;    Blue = 8'h7c;
end 13'he4f:    begin Red = 8'hd5;    Green = 8'h9e;    Blue = 8'h72;
end 13'he50:    begin Red = 8'hdc;    Green = 8'ha2;    Blue = 8'h78;
end 13'he51:    begin Red = 8'hb4;    Green = 8'h9b;    Blue = 8'h78;
end 13'he52:    begin Red = 8'hcf;    Green = 8'haf;    Blue = 8'h84;
end 13'he53:    begin Red = 8'hc7;    Green = 8'ha7;    Blue = 8'h84;
end 13'he54:    begin Red = 8'hab;    Green = 8'h95;    Blue = 8'h6b;
end 13'he55:    begin Red = 8'hc6;    Green = 8'ha5;    Blue = 8'h82;
end 13'he56:    begin Red = 8'h98;    Green = 8'h91;    Blue = 8'h72;
end 13'he57:    begin Red = 8'ha0;    Green = 8'ha3;    Blue = 8'h85;
end 13'he58:    begin Red = 8'h97;    Green = 8'h83;    Blue = 8'h62;
end 13'he59:    begin Red = 8'hb3;    Green = 8'hbf;    Blue = 8'hbf;
end 13'he5a:    begin Red = 8'he6;    Green = 8'hb1;    Blue = 8'h79;
end 13'he5b:    begin Red = 8'h80;    Green = 8'hbb;    Blue = 8'ha3;
end 13'he5c:    begin Red = 8'h92;    Green = 8'hb8;    Blue = 8'h98;
end 13'he5d:    begin Red = 8'he6;    Green = 8'hb9;    Blue = 8'h82;
end 13'he5e:    begin Red = 8'hf1;    Green = 8'hb4;    Blue = 8'h88;
end 13'he5f:    begin Red = 8'hef;    Green = 8'hb3;    Blue = 8'h86;
end 13'he60:    begin Red = 8'hb9;    Green = 8'h84;    Blue = 8'h5d;
end 13'he61:    begin Red = 8'hb3;    Green = 8'h81;    Blue = 8'h56;
end 13'he62:    begin Red = 8'hd3;    Green = 8'he5;    Blue = 8'hc7;
end 13'he63:    begin Red = 8'hd1;    Green = 8'h97;    Blue = 8'h73;
end 13'he64:    begin Red = 8'hc7;    Green = 8'h97;    Blue = 8'h79;
end 13'he65:    begin Red = 8'hd5;    Green = 8'h9b;    Blue = 8'h6d;
end 13'he66:    begin Red = 8'hd8;    Green = 8'h99;    Blue = 8'h6c;
end 13'he67:    begin Red = 8'hb6;    Green = 8'h93;    Blue = 8'h74;
end 13'he68:    begin Red = 8'hd6;    Green = 8'hab;    Blue = 8'h8e;
end 13'he69:    begin Red = 8'hd7;    Green = 8'he2;    Blue = 8'hbf;
end 13'he6a:    begin Red = 8'hdf;    Green = 8'he5;    Blue = 8'hc4;
end 13'he6b:    begin Red = 8'hb5;    Green = 8'h94;    Blue = 8'h6d;
end 13'he6c:    begin Red = 8'hcd;    Green = 8'hac;    Blue = 8'h7b;
end 13'he6d:    begin Red = 8'hdb;    Green = 8'hc6;    Blue = 8'ha3;
end 13'he6e:    begin Red = 8'hcc;    Green = 8'hd6;    Blue = 8'hd2;
end 13'he6f:    begin Red = 8'hdd;    Green = 8'he5;    Blue = 8'hd1;
end 13'he70:    begin Red = 8'hb8;    Green = 8'h8b;    Blue = 8'haf;
end 13'he71:    begin Red = 8'hd0;    Green = 8'h95;    Blue = 8'h6e;
end 13'he72:    begin Red = 8'hd6;    Green = 8'h9b;    Blue = 8'h79;
end 13'he73:    begin Red = 8'hd0;    Green = 8'h9b;    Blue = 8'h75;
end 13'he74:    begin Red = 8'hcf;    Green = 8'h9c;    Blue = 8'h78;
end 13'he75:    begin Red = 8'hd2;    Green = 8'h9b;    Blue = 8'h7b;
end 13'he76:    begin Red = 8'hcf;    Green = 8'ha3;    Blue = 8'h78;
end 13'he77:    begin Red = 8'hd5;    Green = 8'h9e;    Blue = 8'h7d;
end 13'he78:    begin Red = 8'hd3;    Green = 8'ha0;    Blue = 8'h7e;
end 13'he79:    begin Red = 8'hce;    Green = 8'h99;    Blue = 8'h7e;
end 13'he7a:    begin Red = 8'hd2;    Green = 8'ha4;    Blue = 8'h7e;
end 13'he7b:    begin Red = 8'hb1;    Green = 8'h82;    Blue = 8'h5f;
end 13'he7c:    begin Red = 8'ha9;    Green = 8'haf;    Blue = 8'h94;
end 13'he7d:    begin Red = 8'h9d;    Green = 8'hac;    Blue = 8'h93;
end 13'he7e:    begin Red = 8'hef;    Green = 8'hb4;    Blue = 8'h82;
end 13'he7f:    begin Red = 8'hf5;    Green = 8'hb3;    Blue = 8'h85;
end 13'he80:    begin Red = 8'ha4;    Green = 8'h83;    Blue = 8'h5d;
end 13'he81:    begin Red = 8'hb5;    Green = 8'hc7;    Blue = 8'ha7;
end 13'he82:    begin Red = 8'hce;    Green = 8'h9f;    Blue = 8'hc3;
end 13'he83:    begin Red = 8'hbb;    Green = 8'h8e;    Blue = 8'hb0;
end 13'he84:    begin Red = 8'hbd;    Green = 8'h91;    Blue = 8'hb3;
end 13'he85:    begin Red = 8'hd2;    Green = 8'ha4;    Blue = 8'hc8;
end 13'he86:    begin Red = 8'hd2;    Green = 8'ha0;    Blue = 8'hc5;
end 13'he87:    begin Red = 8'ha0;    Green = 8'h7c;    Blue = 8'h96;
end 13'he88:    begin Red = 8'hac;    Green = 8'h86;    Blue = 8'ha7;
end 13'he89:    begin Red = 8'haf;    Green = 8'h85;    Blue = 8'haa;
end 13'he8a:    begin Red = 8'h9d;    Green = 8'h7d;    Blue = 8'h98;
end 13'he8b:    begin Red = 8'hb1;    Green = 8'h8c;    Blue = 8'ha8;
end 13'he8c:    begin Red = 8'hb0;    Green = 8'h8a;    Blue = 8'hac;
end 13'he8d:    begin Red = 8'hd3;    Green = 8'hd4;    Blue = 8'hb4;
end 13'he8e:    begin Red = 8'ha4;    Green = 8'ha8;    Blue = 8'h8f;
end 13'he8f:    begin Red = 8'hc0;    Green = 8'hb4;    Blue = 8'hba;
end 13'he90:    begin Red = 8'hcb;    Green = 8'hd7;    Blue = 8'hd5;
end 13'he91:    begin Red = 8'hb6;    Green = 8'h77;    Blue = 8'h9c;
end 13'he92:    begin Red = 8'hb1;    Green = 8'h78;    Blue = 8'ha8;
end 13'he93:    begin Red = 8'h8f;    Green = 8'h8c;    Blue = 8'h8b;
end 13'he94:    begin Red = 8'hb7;    Green = 8'hab;    Blue = 8'h97;
end 13'he95:    begin Red = 8'h88;    Green = 8'h86;    Blue = 8'h8c;
end 13'he96:    begin Red = 8'h90;    Green = 8'h8c;    Blue = 8'h91;
end 13'he97:    begin Red = 8'h8c;    Green = 8'h8e;    Blue = 8'h85;
end 13'he98:    begin Red = 8'h90;    Green = 8'h8c;    Blue = 8'h98;
end 13'he99:    begin Red = 8'h8a;    Green = 8'h88;    Blue = 8'h8d;
end 13'he9a:    begin Red = 8'h8d;    Green = 8'h8f;    Blue = 8'h8c;
end 13'he9b:    begin Red = 8'hb6;    Green = 8'hac;    Blue = 8'h9c;
end 13'he9c:    begin Red = 8'h8d;    Green = 8'h8b;    Blue = 8'h90;
end 13'he9d:    begin Red = 8'h84;    Green = 8'h8c;    Blue = 8'h8e;
end 13'he9e:    begin Red = 8'hba;    Green = 8'hab;    Blue = 8'h9f;
end 13'he9f:    begin Red = 8'hbb;    Green = 8'had;    Blue = 8'ha3;
end 13'hea0:    begin Red = 8'h8f;    Green = 8'h90;    Blue = 8'h91;
end 13'hea1:    begin Red = 8'h7c;    Green = 8'h7d;    Blue = 8'h7e;
end 13'hea2:    begin Red = 8'h7d;    Green = 8'h80;    Blue = 8'h7c;
end 13'hea3:    begin Red = 8'hc9;    Green = 8'h98;    Blue = 8'h77;
end 13'hea4:    begin Red = 8'h82;    Green = 8'ha6;    Blue = 8'h6f;
end 13'hea5:    begin Red = 8'hc6;    Green = 8'h95;    Blue = 8'hb8;
end 13'hea6:    begin Red = 8'hc1;    Green = 8'h92;    Blue = 8'hb5;
end 13'hea7:    begin Red = 8'hc3;    Green = 8'h95;    Blue = 8'hb6;
end 13'hea8:    begin Red = 8'ha1;    Green = 8'h7b;    Blue = 8'h99;
end 13'hea9:    begin Red = 8'hb2;    Green = 8'h88;    Blue = 8'ha9;
end 13'heaa:    begin Red = 8'hf3;    Green = 8'hdb;    Blue = 8'hb2;
end 13'heab:    begin Red = 8'haf;    Green = 8'h69;    Blue = 8'haa;
end 13'heac:    begin Red = 8'ha9;    Green = 8'h6a;    Blue = 8'h9e;
end 13'head:    begin Red = 8'h7d;    Green = 8'hbf;    Blue = 8'hab;
end 13'heae:    begin Red = 8'hc7;    Green = 8'hb5;    Blue = 8'ha2;
end 13'heaf:    begin Red = 8'h88;    Green = 8'h8b;    Blue = 8'h98;
end 13'heb0:    begin Red = 8'h88;    Green = 8'h8c;    Blue = 8'h89;
end 13'heb1:    begin Red = 8'h90;    Green = 8'h93;    Blue = 8'h97;
end 13'heb2:    begin Red = 8'hcf;    Green = 8'hbc;    Blue = 8'ha7;
end 13'heb3:    begin Red = 8'h89;    Green = 8'h8c;    Blue = 8'h93;
end 13'heb4:    begin Red = 8'h88;    Green = 8'h8f;    Blue = 8'h94;
end 13'heb5:    begin Red = 8'hca;    Green = 8'hbb;    Blue = 8'ha2;
end 13'heb6:    begin Red = 8'hca;    Green = 8'hb6;    Blue = 8'ha6;
end 13'heb7:    begin Red = 8'h8d;    Green = 8'h88;    Blue = 8'h96;
end 13'heb8:    begin Red = 8'h8c;    Green = 8'h94;    Blue = 8'h99;
end 13'heb9:    begin Red = 8'h86;    Green = 8'h90;    Blue = 8'h8e;
end 13'heba:    begin Red = 8'h81;    Green = 8'h89;    Blue = 8'h93;
end 13'hebb:    begin Red = 8'h88;    Green = 8'h8b;    Blue = 8'h8d;
end 13'hebc:    begin Red = 8'h94;    Green = 8'h94;    Blue = 8'h96;
end 13'hebd:    begin Red = 8'h84;    Green = 8'h8e;    Blue = 8'h95;
end 13'hebe:    begin Red = 8'h8e;    Green = 8'h90;    Blue = 8'h9b;
end 13'hebf:    begin Red = 8'hc6;    Green = 8'hbd;    Blue = 8'h98;
end 13'hec0:    begin Red = 8'h7d;    Green = 8'h80;    Blue = 8'h84;
end 13'hec1:    begin Red = 8'h80;    Green = 8'h83;    Blue = 8'h87;
end 13'hec2:    begin Red = 8'h7a;    Green = 8'h82;    Blue = 8'h83;
end 13'hec3:    begin Red = 8'h5c;    Green = 8'h66;    Blue = 8'h50;
end 13'hec4:    begin Red = 8'ha1;    Green = 8'haf;    Blue = 8'h94;
end 13'hec5:    begin Red = 8'h82;    Green = 8'had;    Blue = 8'h7c;
end 13'hec6:    begin Red = 8'h80;    Green = 8'hac;    Blue = 8'h78;
end 13'hec7:    begin Red = 8'h6b;    Green = 8'h92;    Blue = 8'h65;
end 13'hec8:    begin Red = 8'ha9;    Green = 8'h84;    Blue = 8'ha5;
end 13'hec9:    begin Red = 8'h9f;    Green = 8'h78;    Blue = 8'h97;
end 13'heca:    begin Red = 8'had;    Green = 8'h83;    Blue = 8'ha4;
end 13'hecb:    begin Red = 8'hb3;    Green = 8'h84;    Blue = 8'ha8;
end 13'hecc:    begin Red = 8'hbb;    Green = 8'hbf;    Blue = 8'hc9;
end 13'hecd:    begin Red = 8'hb7;    Green = 8'hb4;    Blue = 8'hb3;
end 13'hece:    begin Red = 8'hd8;    Green = 8'hd1;    Blue = 8'hd3;
end 13'hecf:    begin Red = 8'hbb;    Green = 8'h82;    Blue = 8'h57;
end 13'hed0:    begin Red = 8'hb7;    Green = 8'h80;    Blue = 8'h5a;
end 13'hed1:    begin Red = 8'hd3;    Green = 8'h9d;    Blue = 8'h79;
end 13'hed2:    begin Red = 8'hd2;    Green = 8'h9d;    Blue = 8'h6f;
end 13'hed3:    begin Red = 8'h98;    Green = 8'hba;    Blue = 8'h9b;
end 13'hed4:    begin Red = 8'h84;    Green = 8'h69;    Blue = 8'h64;
end 13'hed5:    begin Red = 8'ha6;    Green = 8'h9c;    Blue = 8'h7d;
end 13'hed6:    begin Red = 8'ha9;    Green = 8'h9f;    Blue = 8'h84;
end 13'hed7:    begin Red = 8'h86;    Green = 8'h79;    Blue = 8'h6d;
end 13'hed8:    begin Red = 8'h7d;    Green = 8'h6e;    Blue = 8'h63;
end 13'hed9:    begin Red = 8'h81;    Green = 8'h75;    Blue = 8'h69;
end 13'heda:    begin Red = 8'ha2;    Green = 8'h96;    Blue = 8'h7d;
end 13'hedb:    begin Red = 8'had;    Green = 8'ha2;    Blue = 8'h8b;
end 13'hedc:    begin Red = 8'h7b;    Green = 8'h74;    Blue = 8'h68;
end 13'hedd:    begin Red = 8'h78;    Green = 8'h6d;    Blue = 8'h63;
end 13'hede:    begin Red = 8'h75;    Green = 8'h6a;    Blue = 8'h60;
end 13'hedf:    begin Red = 8'he5;    Green = 8'hbe;    Blue = 8'h8d;
end 13'hee0:    begin Red = 8'hcd;    Green = 8'h94;    Blue = 8'h69;
end 13'hee1:    begin Red = 8'hb2;    Green = 8'h84;    Blue = 8'h65;
end 13'hee2:    begin Red = 8'h75;    Green = 8'h98;    Blue = 8'h6c;
end 13'hee3:    begin Red = 8'hb7;    Green = 8'hc8;    Blue = 8'hae;
end 13'hee4:    begin Red = 8'h6b;    Green = 8'h88;    Blue = 8'h65;
end 13'hee5:    begin Red = 8'hcd;    Green = 8'h9d;    Blue = 8'hc6;
end 13'hee6:    begin Red = 8'h9c;    Green = 8'h79;    Blue = 8'h95;
end 13'hee7:    begin Red = 8'hbb;    Green = 8'hc8;    Blue = 8'hc3;
end 13'hee8:    begin Red = 8'hb3;    Green = 8'h77;    Blue = 8'h9e;
end 13'hee9:    begin Red = 8'haf;    Green = 8'h76;    Blue = 8'h9e;
end 13'heea:    begin Red = 8'h6c;    Green = 8'h63;    Blue = 8'h58;
end 13'heeb:    begin Red = 8'h6c;    Green = 8'h63;    Blue = 8'h5e;
end 13'heec:    begin Red = 8'h91;    Green = 8'hc4;    Blue = 8'haf;
end 13'heed:    begin Red = 8'h8f;    Green = 8'hbb;    Blue = 8'ha3;
end 13'heee:    begin Red = 8'h92;    Green = 8'hb9;    Blue = 8'ha1;
end 13'heef:    begin Red = 8'h97;    Green = 8'hc0;    Blue = 8'ha2;
end 13'hef0:    begin Red = 8'h7e;    Green = 8'h72;    Blue = 8'h70;
end 13'hef1:    begin Red = 8'h87;    Green = 8'h79;    Blue = 8'h73;
end 13'hef2:    begin Red = 8'ha7;    Green = 8'ha0;    Blue = 8'h7c;
end 13'hef3:    begin Red = 8'h79;    Green = 8'h69;    Blue = 8'h62;
end 13'hef4:    begin Red = 8'hd8;    Green = 8'ha3;    Blue = 8'h78;
end 13'hef5:    begin Red = 8'hc7;    Green = 8'hac;    Blue = 8'h82;
end 13'hef6:    begin Red = 8'h86;    Green = 8'h93;    Blue = 8'h74;
end 13'hef7:    begin Red = 8'ha3;    Green = 8'h80;    Blue = 8'h69;
end 13'hef8:    begin Red = 8'hb9;    Green = 8'hc3;    Blue = 8'h9e;
end 13'hef9:    begin Red = 8'h97;    Green = 8'h9a;    Blue = 8'h72;
end 13'hefa:    begin Red = 8'ha9;    Green = 8'h82;    Blue = 8'h6a;
end 13'hefb:    begin Red = 8'hc9;    Green = 8'h92;    Blue = 8'h78;
end 13'hefc:    begin Red = 8'hce;    Green = 8'h94;    Blue = 8'h71;
end 13'hefd:    begin Red = 8'h8c;    Green = 8'hb3;    Blue = 8'h87;
end 13'hefe:    begin Red = 8'hd0;    Green = 8'ha1;    Blue = 8'hc7;
end 13'heff:    begin Red = 8'hc1;    Green = 8'hbf;    Blue = 8'hca;
end 13'hf00:    begin Red = 8'hbb;    Green = 8'h84;    Blue = 8'hac;
end 13'hf01:    begin Red = 8'hb6;    Green = 8'h82;    Blue = 8'hb5;
end 13'hf02:    begin Red = 8'hdd;    Green = 8'he5;    Blue = 8'he1;
end 13'hf03:    begin Red = 8'ha1;    Green = 8'hc5;    Blue = 8'hac;
end 13'hf04:    begin Red = 8'hab;    Green = 8'ha3;    Blue = 8'h87;
end 13'hf05:    begin Red = 8'h7a;    Green = 8'h69;    Blue = 8'h5e;
end 13'hf06:    begin Red = 8'hdc;    Green = 8'ha0;    Blue = 8'h87;
end 13'hf07:    begin Red = 8'hca;    Green = 8'had;    Blue = 8'h81;
end 13'hf08:    begin Red = 8'h85;    Green = 8'h91;    Blue = 8'h78;
end 13'hf09:    begin Red = 8'hc7;    Green = 8'h99;    Blue = 8'h75;
end 13'hf0a:    begin Red = 8'haf;    Green = 8'h88;    Blue = 8'h6e;
end 13'hf0b:    begin Red = 8'hbb;    Green = 8'hd6;    Blue = 8'hb9;
end 13'hf0c:    begin Red = 8'h94;    Green = 8'ha1;    Blue = 8'h88;
end 13'hf0d:    begin Red = 8'hae;    Green = 8'h86;    Blue = 8'h6a;
end 13'hf0e:    begin Red = 8'hc5;    Green = 8'h98;    Blue = 8'h70;
end 13'hf0f:    begin Red = 8'hab;    Green = 8'h7a;    Blue = 8'h9b;
end 13'hf10:    begin Red = 8'ha4;    Green = 8'h5b;    Blue = 8'h90;
end 13'hf11:    begin Red = 8'hc8;    Green = 8'hb0;    Blue = 8'h88;
end 13'hf12:    begin Red = 8'hc1;    Green = 8'hb1;    Blue = 8'h89;
end 13'hf13:    begin Red = 8'haa;    Green = 8'h97;    Blue = 8'h7c;
end 13'hf14:    begin Red = 8'hab;    Green = 8'haa;    Blue = 8'h85;
end 13'hf15:    begin Red = 8'h8d;    Green = 8'h90;    Blue = 8'h7d;
end 13'hf16:    begin Red = 8'he5;    Green = 8'hf0;    Blue = 8'hc6;
end 13'hf17:    begin Red = 8'hb5;    Green = 8'hbd;    Blue = 8'ha0;
end 13'hf18:    begin Red = 8'h84;    Green = 8'h76;    Blue = 8'h6c;
end 13'hf19:    begin Red = 8'he9;    Green = 8'he4;    Blue = 8'hbe;
end 13'hf1a:    begin Red = 8'hbe;    Green = 8'hb8;    Blue = 8'h99;
end 13'hf1b:    begin Red = 8'h7d;    Green = 8'h76;    Blue = 8'h6f;
end 13'hf1c:    begin Red = 8'h8c;    Green = 8'hab;    Blue = 8'he3;
end 13'hf1d:    begin Red = 8'ha9;    Green = 8'h9a;    Blue = 8'h7a;
end 13'hf1e:    begin Red = 8'hbe;    Green = 8'hc3;    Blue = 8'hcf;
end 13'hf1f:    begin Red = 8'hc7;    Green = 8'hd1;    Blue = 8'hc6;
end 13'hf20:    begin Red = 8'hc0;    Green = 8'hcf;    Blue = 8'hbe;
end 13'hf21:    begin Red = 8'had;    Green = 8'h71;    Blue = 8'h9f;
end 13'hf22:    begin Red = 8'had;    Green = 8'h5f;    Blue = 8'h8e;
end 13'hf23:    begin Red = 8'h9d;    Green = 8'hc2;    Blue = 8'ha5;
end 13'hf24:    begin Red = 8'h8f;    Green = 8'hbd;    Blue = 8'h94;
end 13'hf25:    begin Red = 8'hf1;    Green = 8'he9;    Blue = 8'hd5;
end 13'hf26:    begin Red = 8'hd3;    Green = 8'hce;    Blue = 8'hbb;
end 13'hf27:    begin Red = 8'hd6;    Green = 8'hd2;    Blue = 8'hc0;
end 13'hf28:    begin Red = 8'hd6;    Green = 8'hcf;    Blue = 8'hbd;
end 13'hf29:    begin Red = 8'hb1;    Green = 8'ha7;    Blue = 8'h98;
end 13'hf2a:    begin Red = 8'hac;    Green = 8'had;    Blue = 8'h94;
end 13'hf2b:    begin Red = 8'hce;    Green = 8'hbd;    Blue = 8'h95;
end 13'hf2c:    begin Red = 8'hb1;    Green = 8'ha5;    Blue = 8'h84;
end 13'hf2d:    begin Red = 8'hdf;    Green = 8'he5;    Blue = 8'hbb;
end 13'hf2e:    begin Red = 8'haf;    Green = 8'h81;    Blue = 8'h6a;
end 13'hf2f:    begin Red = 8'h71;    Green = 8'h73;    Blue = 8'h64;
end 13'hf30:    begin Red = 8'hdf;    Green = 8'hd9;    Blue = 8'hb2;
end 13'hf31:    begin Red = 8'he3;    Green = 8'hdc;    Blue = 8'hbb;
end 13'hf32:    begin Red = 8'hba;    Green = 8'hb4;    Blue = 8'h91;
end 13'hf33:    begin Red = 8'hbd;    Green = 8'ha7;    Blue = 8'h85;
end 13'hf34:    begin Red = 8'hb4;    Green = 8'ha7;    Blue = 8'h84;
end 13'hf35:    begin Red = 8'hc3;    Green = 8'hc4;    Blue = 8'hd0;
end 13'hf36:    begin Red = 8'hbe;    Green = 8'hb6;    Blue = 8'hb9;
end 13'hf37:    begin Red = 8'hbb;    Green = 8'h88;    Blue = 8'hb3;
end 13'hf38:    begin Red = 8'hb7;    Green = 8'h83;    Blue = 8'h9e;
end 13'hf39:    begin Red = 8'haa;    Green = 8'h76;    Blue = 8'ha3;
end 13'hf3a:    begin Red = 8'ha2;    Green = 8'h88;    Blue = 8'h6f;
end 13'hf3b:    begin Red = 8'hf2;    Green = 8'he1;    Blue = 8'hce;
end 13'hf3c:    begin Red = 8'he2;    Green = 8'hd8;    Blue = 8'hc3;
end 13'hf3d:    begin Red = 8'hcf;    Green = 8'hc6;    Blue = 8'hb1;
end 13'hf3e:    begin Red = 8'hd2;    Green = 8'hc9;    Blue = 8'hb4;
end 13'hf3f:    begin Red = 8'had;    Green = 8'ha6;    Blue = 8'h98;
end 13'hf40:    begin Red = 8'hae;    Green = 8'ha5;    Blue = 8'h95;
end 13'hf41:    begin Red = 8'had;    Green = 8'haf;    Blue = 8'h97;
end 13'hf42:    begin Red = 8'hc4;    Green = 8'hb3;    Blue = 8'h8e;
end 13'hf43:    begin Red = 8'ha8;    Green = 8'haf;    Blue = 8'h98;
end 13'hf44:    begin Red = 8'ha7;    Green = 8'h8e;    Blue = 8'h61;
end 13'hf45:    begin Red = 8'hb3;    Green = 8'h99;    Blue = 8'h7a;
end 13'hf46:    begin Red = 8'hbb;    Green = 8'hb5;    Blue = 8'h94;
end 13'hf47:    begin Red = 8'h6b;    Green = 8'h78;    Blue = 8'h9f;
end 13'hf48:    begin Red = 8'h68;    Green = 8'h7f;    Blue = 8'h9f;
end 13'hf49:    begin Red = 8'h91;    Green = 8'hb6;    Blue = 8'hf3;
end 13'hf4a:    begin Red = 8'h8c;    Green = 8'ha8;    Blue = 8'he6;
end 13'hf4b:    begin Red = 8'h95;    Green = 8'h71;    Blue = 8'h94;
end 13'hf4c:    begin Red = 8'h96;    Green = 8'h71;    Blue = 8'h8e;
end 13'hf4d:    begin Red = 8'h8a;    Green = 8'h65;    Blue = 8'h82;
end 13'hf4e:    begin Red = 8'h8c;    Green = 8'h69;    Blue = 8'h84;
end 13'hf4f:    begin Red = 8'h87;    Green = 8'h6f;    Blue = 8'h84;
end 13'hf50:    begin Red = 8'h90;    Green = 8'h71;    Blue = 8'h8e;
end 13'hf51:    begin Red = 8'h94;    Green = 8'h6f;    Blue = 8'h8c;
end 13'hf52:    begin Red = 8'h93;    Green = 8'h6c;    Blue = 8'h8b;
end 13'hf53:    begin Red = 8'h98;    Green = 8'h6e;    Blue = 8'h91;
end 13'hf54:    begin Red = 8'hde;    Green = 8'hd1;    Blue = 8'ha7;
end 13'hf55:    begin Red = 8'h85;    Green = 8'h75;    Blue = 8'h74;
end 13'hf56:    begin Red = 8'h62;    Green = 8'h7d;    Blue = 8'h9b;
end 13'hf57:    begin Red = 8'h90;    Green = 8'hac;    Blue = 8'hf9;
end 13'hf58:    begin Red = 8'h8e;    Green = 8'had;    Blue = 8'hec;
end 13'hf59:    begin Red = 8'h9b;    Green = 8'h85;    Blue = 8'h61;
end 13'hf5a:    begin Red = 8'hda;    Green = 8'he7;    Blue = 8'he7;
end 13'hf5b:    begin Red = 8'h8f;    Green = 8'h88;    Blue = 8'h80;
end 13'hf5c:    begin Red = 8'hcd;    Green = 8'hc7;    Blue = 8'hb3;
end 13'hf5d:    begin Red = 8'hff;    Green = 8'hf3;    Blue = 8'hdc;
end 13'hf5e:    begin Red = 8'hf2;    Green = 8'he7;    Blue = 8'hd0;
end 13'hf5f:    begin Red = 8'h9e;    Green = 8'h92;    Blue = 8'h80;
end 13'hf60:    begin Red = 8'he8;    Green = 8'hdf;    Blue = 8'hc9;
end 13'hf61:    begin Red = 8'he3;    Green = 8'hdf;    Blue = 8'hc8;
end 13'hf62:    begin Red = 8'hbf;    Green = 8'hb8;    Blue = 8'hab;
end 13'hf63:    begin Red = 8'hc7;    Green = 8'hc0;    Blue = 8'hae;
end 13'hf64:    begin Red = 8'hbe;    Green = 8'hb8;    Blue = 8'ha6;
end 13'hf65:    begin Red = 8'hf1;    Green = 8'hee;    Blue = 8'hd9;
end 13'hf66:    begin Red = 8'h5a;    Green = 8'h78;    Blue = 8'ha3;
end 13'hf67:    begin Red = 8'h94;    Green = 8'hba;    Blue = 8'hff;
end 13'hf68:    begin Red = 8'h8c;    Green = 8'haf;    Blue = 8'hfa;
end 13'hf69:    begin Red = 8'h90;    Green = 8'hb3;    Blue = 8'hff;
end 13'hf6a:    begin Red = 8'h9b;    Green = 8'h82;    Blue = 8'h71;
end 13'hf6b:    begin Red = 8'h85;    Green = 8'h5d;    Blue = 8'h90;
end 13'hf6c:    begin Red = 8'h82;    Green = 8'h5a;    Blue = 8'h87;
end 13'hf6d:    begin Red = 8'h79;    Green = 8'h52;    Blue = 8'h7f;
end 13'hf6e:    begin Red = 8'h7c;    Green = 8'h4e;    Blue = 8'h7a;
end 13'hf6f:    begin Red = 8'h8b;    Green = 8'h5f;    Blue = 8'h93;
end 13'hf70:    begin Red = 8'h8c;    Green = 8'h61;    Blue = 8'h8c;
end 13'hf71:    begin Red = 8'h89;    Green = 8'h5d;    Blue = 8'h89;
end 13'hf72:    begin Red = 8'h80;    Green = 8'h58;    Blue = 8'h82;
end 13'hf73:    begin Red = 8'h81;    Green = 8'h55;    Blue = 8'h81;
end 13'hf74:    begin Red = 8'h8a;    Green = 8'h5e;    Blue = 8'h8c;
end 13'hf75:    begin Red = 8'h8f;    Green = 8'h5e;    Blue = 8'h94;
end 13'hf76:    begin Red = 8'he5;    Green = 8'hcf;    Blue = 8'ha9;
end 13'hf77:    begin Red = 8'h59;    Green = 8'h74;    Blue = 8'ha6;
end 13'hf78:    begin Red = 8'h95;    Green = 8'hbc;    Blue = 8'hfb;
end 13'hf79:    begin Red = 8'h93;    Green = 8'had;    Blue = 8'hff;
end 13'hf7a:    begin Red = 8'hc5;    Green = 8'hd3;    Blue = 8'hc7;
end 13'hf7b:    begin Red = 8'hc1;    Green = 8'hcb;    Blue = 8'hc4;
end 13'hf7c:    begin Red = 8'hd9;    Green = 8'he6;    Blue = 8'hde;
end 13'hf7d:    begin Red = 8'h80;    Green = 8'h7c;    Blue = 8'h6a;
end 13'hf7e:    begin Red = 8'hb3;    Green = 8'hab;    Blue = 8'h99;
end 13'hf7f:    begin Red = 8'hc9;    Green = 8'hbf;    Blue = 8'hab;
end 13'hf80:    begin Red = 8'hd4;    Green = 8'hca;    Blue = 8'hb6;
end 13'hf81:    begin Red = 8'ha9;    Green = 8'h9c;    Blue = 8'h90;
end 13'hf82:    begin Red = 8'ha9;    Green = 8'h9c;    Blue = 8'h88;
end 13'hf83:    begin Red = 8'hb3;    Green = 8'hb3;    Blue = 8'h98;
end 13'hf84:    begin Red = 8'heb;    Green = 8'he2;    Blue = 8'hcc;
end 13'hf85:    begin Red = 8'hed;    Green = 8'he4;    Blue = 8'hce;
end 13'hf86:    begin Red = 8'hcc;    Green = 8'hc4;    Blue = 8'hb0;
end 13'hf87:    begin Red = 8'hea;    Green = 8'he9;    Blue = 8'hb3;
end 13'hf88:    begin Red = 8'hdf;    Green = 8'hc7;    Blue = 8'h9c;
end 13'hf89:    begin Red = 8'hdd;    Green = 8'hc5;    Blue = 8'h9d;
end 13'hf8a:    begin Red = 8'hea;    Green = 8'hca;    Blue = 8'ha5;
end 13'hf8b:    begin Red = 8'hbf;    Green = 8'haf;    Blue = 8'h98;
end 13'hf8c:    begin Red = 8'hd6;    Green = 8'hd7;    Blue = 8'hb2;
end 13'hf8d:    begin Red = 8'h7d;    Green = 8'h75;    Blue = 8'h74;
end 13'hf8e:    begin Red = 8'ha4;    Green = 8'h76;    Blue = 8'h94;
end 13'hf8f:    begin Red = 8'ha0;    Green = 8'h6f;    Blue = 8'h96;
end 13'hf90:    begin Red = 8'hb5;    Green = 8'h82;    Blue = 8'haa;
end 13'hf91:    begin Red = 8'haf;    Green = 8'h6f;    Blue = 8'h99;
end 13'hf92:    begin Red = 8'hd7;    Green = 8'hcc;    Blue = 8'hb7;
end 13'hf93:    begin Red = 8'hd5;    Green = 8'hcc;    Blue = 8'hbc;
end 13'hf94:    begin Red = 8'hba;    Green = 8'haf;    Blue = 8'ha0;
end 13'hf95:    begin Red = 8'he4;    Green = 8'hdd;    Blue = 8'hc6;
end 13'hf96:    begin Red = 8'h6b;    Green = 8'h60;    Blue = 8'h59;
end 13'hf97:    begin Red = 8'hce;    Green = 8'hc2;    Blue = 8'ha7;
end 13'hf98:    begin Red = 8'hca;    Green = 8'hbe;    Blue = 8'ha7;
end 13'hf99:    begin Red = 8'ha2;    Green = 8'ha7;    Blue = 8'h87;
end 13'hf9a:    begin Red = 8'h47;    Green = 8'h40;    Blue = 8'h44;
end 13'hf9b:    begin Red = 8'hb4;    Green = 8'haf;    Blue = 8'h8d;
end 13'hf9c:    begin Red = 8'h61;    Green = 8'h77;    Blue = 8'h94;
end 13'hf9d:    begin Red = 8'hf0;    Green = 8'hdb;    Blue = 8'hb4;
end 13'hf9e:    begin Red = 8'hbb;    Green = 8'hae;    Blue = 8'h85;
end 13'hf9f:    begin Red = 8'h9b;    Green = 8'ha2;    Blue = 8'hae;
end 13'hfa0:    begin Red = 8'ha9;    Green = 8'ha7;    Blue = 8'hb0;
end 13'hfa1:    begin Red = 8'hb0;    Green = 8'ha5;    Blue = 8'hb1;
end 13'hfa2:    begin Red = 8'hee;    Green = 8'he6;    Blue = 8'hd2;
end 13'hfa3:    begin Red = 8'hf0;    Green = 8'he5;    Blue = 8'hd6;
end 13'hfa4:    begin Red = 8'hf5;    Green = 8'hec;    Blue = 8'hd6;
end 13'hfa5:    begin Red = 8'hb8;    Green = 8'haf;    Blue = 8'h9d;
end 13'hfa6:    begin Red = 8'hee;    Green = 8'he8;    Blue = 8'hd7;
end 13'hfa7:    begin Red = 8'he5;    Green = 8'hdd;    Blue = 8'hc1;
end 13'hfa8:    begin Red = 8'he2;    Green = 8'he1;    Blue = 8'hca;
end 13'hfa9:    begin Red = 8'he3;    Green = 8'hdc;    Blue = 8'hce;
end 13'hfaa:    begin Red = 8'hf5;    Green = 8'hf4;    Blue = 8'he3;
end 13'hfab:    begin Red = 8'h88;    Green = 8'ha5;    Blue = 8'h8c;
end 13'hfac:    begin Red = 8'h8c;    Green = 8'h90;    Blue = 8'h8f;
end 13'hfad:    begin Red = 8'hb6;    Green = 8'hb6;    Blue = 8'h99;
end 13'hfae:    begin Red = 8'hc0;    Green = 8'hb7;    Blue = 8'ha0;
end 13'hfaf:    begin Red = 8'hca;    Green = 8'hbf;    Blue = 8'hb3;
end 13'hfb0:    begin Red = 8'h75;    Green = 8'h60;    Blue = 8'h51;
end 13'hfb1:    begin Red = 8'hd1;    Green = 8'hdd;    Blue = 8'hc3;
end 13'hfb2:    begin Red = 8'h79;    Green = 8'h65;    Blue = 8'h57;
end 13'hfb3:    begin Red = 8'h98;    Green = 8'h8d;    Blue = 8'h71;
end 13'hfb4:    begin Red = 8'ha2;    Green = 8'h9c;    Blue = 8'h86;
end 13'hfb5:    begin Red = 8'h58;    Green = 8'h79;    Blue = 8'ha9;
end 13'hfb6:    begin Red = 8'hc3;    Green = 8'had;    Blue = 8'h85;
end 13'hfb7:    begin Red = 8'hac;    Green = 8'h95;    Blue = 8'h72;
end 13'hfb8:    begin Red = 8'hb5;    Green = 8'h98;    Blue = 8'h82;
end 13'hfb9:    begin Red = 8'heb;    Green = 8'hde;    Blue = 8'had;
end 13'hfba:    begin Red = 8'h62;    Green = 8'h71;    Blue = 8'ha0;
end 13'hfbb:    begin Red = 8'ha5;    Green = 8'h88;    Blue = 8'h78;
end 13'hfbc:    begin Red = 8'ha0;    Green = 8'ha3;    Blue = 8'ha8;
end 13'hfbd:    begin Red = 8'hff;    Green = 8'hf9;    Blue = 8'hf1;
end 13'hfbe:    begin Red = 8'hfd;    Green = 8'hf8;    Blue = 8'hed;
end 13'hfbf:    begin Red = 8'hf0;    Green = 8'he5;    Blue = 8'hca;
end 13'hfc0:    begin Red = 8'hfc;    Green = 8'hf6;    Blue = 8'he5;
end 13'hfc1:    begin Red = 8'hfc;    Green = 8'hfb;    Blue = 8'he5;
end 13'hfc2:    begin Red = 8'hf7;    Green = 8'hed;    Blue = 8'hda;
end 13'hfc3:    begin Red = 8'hf5;    Green = 8'hea;    Blue = 8'hdd;
end 13'hfc4:    begin Red = 8'he5;    Green = 8'hde;    Blue = 8'hd0;
end 13'hfc5:    begin Red = 8'he8;    Green = 8'he1;    Blue = 8'hd2;
end 13'hfc6:    begin Red = 8'he1;    Green = 8'hde;    Blue = 8'hcf;
end 13'hfc7:    begin Red = 8'hff;    Green = 8'hfb;    Blue = 8'hec;
end 13'hfc8:    begin Red = 8'hf9;    Green = 8'hf3;    Blue = 8'he2;
end 13'hfc9:    begin Red = 8'h96;    Green = 8'h99;    Blue = 8'ha0;
end 13'hfca:    begin Red = 8'h98;    Green = 8'h9c;    Blue = 8'h9c;
end 13'hfcb:    begin Red = 8'h96;    Green = 8'h99;    Blue = 8'h9a;
end 13'hfcc:    begin Red = 8'h94;    Green = 8'h97;    Blue = 8'h99;
end 13'hfcd:    begin Red = 8'hb3;    Green = 8'hb4;    Blue = 8'h94;
end 13'hfce:    begin Red = 8'h93;    Green = 8'h98;    Blue = 8'h80;
end 13'hfcf:    begin Red = 8'hc6;    Green = 8'hbd;    Blue = 8'ha5;
end 13'hfd0:    begin Red = 8'hcc;    Green = 8'hc9;    Blue = 8'hb5;
end 13'hfd1:    begin Red = 8'hbf;    Green = 8'hc9;    Blue = 8'ha3;
end 13'hfd2:    begin Red = 8'ha1;    Green = 8'haa;    Blue = 8'h8a;
end 13'hfd3:    begin Red = 8'hf3;    Green = 8'hf0;    Blue = 8'hda;
end 13'hfd4:    begin Red = 8'hde;    Green = 8'hb4;    Blue = 8'h8f;
end 13'hfd5:    begin Red = 8'h7d;    Green = 8'h67;    Blue = 8'h56;
end 13'hfd6:    begin Red = 8'hd5;    Green = 8'he1;    Blue = 8'hc7;
end 13'hfd7:    begin Red = 8'ha6;    Green = 8'h87;    Blue = 8'h68;
end 13'hfd8:    begin Red = 8'h7c;    Green = 8'h6e;    Blue = 8'h68;
end 13'hfd9:    begin Red = 8'hf3;    Green = 8'hd4;    Blue = 8'hb3;
end 13'hfda:    begin Red = 8'hae;    Green = 8'ha7;    Blue = 8'h9d;
end 13'hfdb:    begin Red = 8'hb7;    Green = 8'haa;    Blue = 8'ha0;
end 13'hfdc:    begin Red = 8'hb7;    Green = 8'ha8;    Blue = 8'ha3;
end 13'hfdd:    begin Red = 8'hf0;    Green = 8'hd6;    Blue = 8'haf;
end 13'hfde:    begin Red = 8'hb3;    Green = 8'hb8;    Blue = 8'hc2;
end 13'hfdf:    begin Red = 8'hf3;    Green = 8'he2;    Blue = 8'hd5;
end 13'hfe0:    begin Red = 8'hed;    Green = 8'he9;    Blue = 8'hd4;
end 13'hfe1:    begin Red = 8'ha1;    Green = 8'h8c;    Blue = 8'h60;
end 13'hfe2:    begin Red = 8'h9e;    Green = 8'h8c;    Blue = 8'h65;
end 13'hfe3:    begin Red = 8'h8b;    Green = 8'h7b;    Blue = 8'h44;
end 13'hfe4:    begin Red = 8'hff;    Green = 8'hfd;    Blue = 8'hf0;
end 13'hfe5:    begin Red = 8'he6;    Green = 8'hdd;    Blue = 8'hca;
end 13'hfe6:    begin Red = 8'hdd;    Green = 8'hd1;    Blue = 8'h9b;
end 13'hfe7:    begin Red = 8'he0;    Green = 8'hcf;    Blue = 8'h9d;
end 13'hfe8:    begin Red = 8'hdf;    Green = 8'hcb;    Blue = 8'h98;
end 13'hfe9:    begin Red = 8'h4e;    Green = 8'h43;    Blue = 8'h41;
end 13'hfea:    begin Red = 8'h5a;    Green = 8'h52;    Blue = 8'h4e;
end 13'hfeb:    begin Red = 8'h99;    Green = 8'h73;    Blue = 8'h55;
end 13'hfec:    begin Red = 8'hd1;    Green = 8'hb2;    Blue = 8'h91;
end 13'hfed:    begin Red = 8'hd8;    Green = 8'hc0;    Blue = 8'h98;
end 13'hfee:    begin Red = 8'hc1;    Green = 8'hb9;    Blue = 8'haf;
end 13'hfef:    begin Red = 8'hc3;    Green = 8'hbb;    Blue = 8'hb3;
end 13'hff0:    begin Red = 8'hc7;    Green = 8'hbb;    Blue = 8'hbb;
end 13'hff1:    begin Red = 8'hbf;    Green = 8'h95;    Blue = 8'h7a;
end 13'hff2:    begin Red = 8'hbf;    Green = 8'h90;    Blue = 8'h60;
end 13'hff3:    begin Red = 8'hb3;    Green = 8'h9e;    Blue = 8'h77;
end 13'hff4:    begin Red = 8'hf1;    Green = 8'hd2;    Blue = 8'hb8;
end 13'hff5:    begin Red = 8'he9;    Green = 8'hce;    Blue = 8'hae;
end 13'hff6:    begin Red = 8'hb3;    Green = 8'hba;    Blue = 8'hbb;
end 13'hff7:    begin Red = 8'hb3;    Green = 8'hb0;    Blue = 8'hb1;
end 13'hff8:    begin Red = 8'h8d;    Green = 8'h7d;    Blue = 8'h3e;
end 13'hff9:    begin Red = 8'h7f;    Green = 8'h61;    Blue = 8'h3a;
end 13'hffa:    begin Red = 8'hf5;    Green = 8'he7;    Blue = 8'hd7;
end 13'hffb:    begin Red = 8'hea;    Green = 8'he3;    Blue = 8'hd5;
end 13'hffc:    begin Red = 8'h90;    Green = 8'h7e;    Blue = 8'h44;
end 13'hffd:    begin Red = 8'h89;    Green = 8'h6c;    Blue = 8'h3f;
end 13'hffe:    begin Red = 8'hef;    Green = 8'hea;    Blue = 8'hdd;
end 13'hfff:    begin Red = 8'he8;    Green = 8'hdf;    Blue = 8'hce;
end 13'h1000:    begin Red = 8'he4;    Green = 8'hd9;    Blue = 8'hcc;
end 13'h1001:    begin Red = 8'hc1;    Green = 8'hb7;    Blue = 8'ha4;
end 13'h1002:    begin Red = 8'ha7;    Green = 8'ha7;    Blue = 8'h8e;
end 13'h1003:    begin Red = 8'ha9;    Green = 8'h87;    Blue = 8'h63;
end 13'h1004:    begin Red = 8'hdf;    Green = 8'he0;    Blue = 8'hc0;
end 13'h1005:    begin Red = 8'hb1;    Green = 8'ha9;    Blue = 8'ha1;
end 13'h1006:    begin Red = 8'haf;    Green = 8'ha9;    Blue = 8'ha7;
end 13'h1007:    begin Red = 8'hc6;    Green = 8'hb8;    Blue = 8'hb2;
end 13'h1008:    begin Red = 8'hb5;    Green = 8'ha3;    Blue = 8'h7b;
end 13'h1009:    begin Red = 8'hbc;    Green = 8'h97;    Blue = 8'h6d;
end 13'h100a:    begin Red = 8'hc3;    Green = 8'hb9;    Blue = 8'hac;
end 13'h100b:    begin Red = 8'hc0;    Green = 8'hbc;    Blue = 8'had;
end 13'h100c:    begin Red = 8'h9d;    Green = 8'h9e;    Blue = 8'hae;
end 13'h100d:    begin Red = 8'ha5;    Green = 8'ha6;    Blue = 8'haa;
end 13'h100e:    begin Red = 8'hc6;    Green = 8'hb9;    Blue = 8'hc1;
end 13'h100f:    begin Red = 8'h98;    Green = 8'h8c;    Blue = 8'h61;
end 13'h1010:    begin Red = 8'ha1;    Green = 8'h89;    Blue = 8'h5e;
end 13'h1011:    begin Red = 8'h99;    Green = 8'h8b;    Blue = 8'h66;
end 13'h1012:    begin Red = 8'h88;    Green = 8'h78;    Blue = 8'h42;
end 13'h1013:    begin Red = 8'h9e;    Green = 8'h8f;    Blue = 8'h62;
end 13'h1014:    begin Red = 8'hba;    Green = 8'hb0;    Blue = 8'h9b;
end 13'h1015:    begin Red = 8'hfe;    Green = 8'hf7;    Blue = 8'he9;
end 13'h1016:    begin Red = 8'h80;    Green = 8'ha8;    Blue = 8'h8a;
end 13'h1017:    begin Red = 8'h9d;    Green = 8'h92;    Blue = 8'h7b;
end 13'h1018:    begin Red = 8'h48;    Green = 8'h47;    Blue = 8'h44;
end 13'h1019:    begin Red = 8'hbe;    Green = 8'hc9;    Blue = 8'h9f;
end 13'h101a:    begin Red = 8'hc4;    Green = 8'hb4;    Blue = 8'hac;
end 13'h101b:    begin Red = 8'hb7;    Green = 8'hbd;    Blue = 8'hac;
end 13'h101c:    begin Red = 8'hca;    Green = 8'hce;    Blue = 8'hc0;
end 13'h101d:    begin Red = 8'hd6;    Green = 8'hc5;    Blue = 8'hbb;
end 13'h101e:    begin Red = 8'hce;    Green = 8'hcd;    Blue = 8'hbc;
end 13'h101f:    begin Red = 8'hd3;    Green = 8'hc7;    Blue = 8'hc5;
end 13'h1020:    begin Red = 8'hbc;    Green = 8'h9f;    Blue = 8'h7c;
end 13'h1021:    begin Red = 8'hde;    Green = 8'hd1;    Blue = 8'hc7;
end 13'h1022:    begin Red = 8'hd0;    Green = 8'hc7;    Blue = 8'hbb;
end 13'h1023:    begin Red = 8'hf5;    Green = 8'hec;    Blue = 8'hc8;
end 13'h1024:    begin Red = 8'ha0;    Green = 8'h8c;    Blue = 8'h5b;
end 13'h1025:    begin Red = 8'hf1;    Green = 8'he3;    Blue = 8'hdb;
end 13'h1026:    begin Red = 8'hfc;    Green = 8'hfc;    Blue = 8'hf6;
end 13'h1027:    begin Red = 8'hf7;    Green = 8'hf4;    Blue = 8'he0;
end 13'h1028:    begin Red = 8'hfa;    Green = 8'hf6;    Blue = 8'he1;
end 13'h1029:    begin Red = 8'h98;    Green = 8'h9b;    Blue = 8'h7d;
end 13'h102a:    begin Red = 8'hba;    Green = 8'hc4;    Blue = 8'hae;
end 13'h102b:    begin Red = 8'haf;    Green = 8'h8c;    Blue = 8'h54;
end 13'h102c:    begin Red = 8'hcd;    Green = 8'hcb;    Blue = 8'hc1;
end 13'h102d:    begin Red = 8'hab;    Green = 8'hb3;    Blue = 8'hba;
end 13'h102e:    begin Red = 8'hb2;    Green = 8'hb3;    Blue = 8'hbd;
end 13'h102f:    begin Red = 8'hae;    Green = 8'haf;    Blue = 8'hb9;
end 13'h1030:    begin Red = 8'hd2;    Green = 8'hd4;    Blue = 8'hde;
end 13'h1031:    begin Red = 8'hc7;    Green = 8'hca;    Blue = 8'he0;
end 13'h1032:    begin Red = 8'hef;    Green = 8'he2;    Blue = 8'hd3;
end 13'h1033:    begin Red = 8'h8a;    Green = 8'h76;    Blue = 8'h41;
end 13'h1034:    begin Red = 8'hfe;    Green = 8'hf2;    Blue = 8'hed;
end 13'h1035:    begin Red = 8'hff;    Green = 8'hff;    Blue = 8'hf3;
end 13'h1036:    begin Red = 8'h90;    Green = 8'h98;    Blue = 8'h99;
end 13'h1037:    begin Red = 8'hc9;    Green = 8'hb7;    Blue = 8'h8f;
end 13'h1038:    begin Red = 8'hbf;    Green = 8'h9c;    Blue = 8'h78;
end 13'h1039:    begin Red = 8'hd3;    Green = 8'hc9;    Blue = 8'hbb;
end 13'h103a:    begin Red = 8'hd1;    Green = 8'hc9;    Blue = 8'hac;
end 13'h103b:    begin Red = 8'hd3;    Green = 8'hc9;    Blue = 8'hc2;
end 13'h103c:    begin Red = 8'hf5;    Green = 8'hf0;    Blue = 8'he6;
end 13'h103d:    begin Red = 8'he8;    Green = 8'hd9;    Blue = 8'hcb;
end 13'h103e:    begin Red = 8'hd3;    Green = 8'hc4;    Blue = 8'hb7;
end 13'h103f:    begin Red = 8'he4;    Green = 8'he2;    Blue = 8'hc7;
end 13'h1040:    begin Red = 8'he2;    Green = 8'he4;    Blue = 8'hc0;
end 13'h1041:    begin Red = 8'h8a;    Green = 8'h75;    Blue = 8'h5d;
end 13'h1042:    begin Red = 8'hb8;    Green = 8'hb4;    Blue = 8'haf;
end 13'h1043:    begin Red = 8'hdf;    Green = 8'hc0;    Blue = 8'h93;
end 13'h1044:    begin Red = 8'h7f;    Green = 8'h69;    Blue = 8'h52;
end 13'h1045:    begin Red = 8'hea;    Green = 8'hd5;    Blue = 8'ha9;
end 13'h1046:    begin Red = 8'hf1;    Green = 8'hd5;    Blue = 8'ha8;
end 13'h1047:    begin Red = 8'hf4;    Green = 8'hd6;    Blue = 8'hac;
end 13'h1048:    begin Red = 8'he5;    Green = 8'hca;    Blue = 8'ha0;
end 13'h1049:    begin Red = 8'hdb;    Green = 8'hbb;    Blue = 8'h91;
end 13'h104a:    begin Red = 8'hda;    Green = 8'hbe;    Blue = 8'h94;
end 13'h104b:    begin Red = 8'h92;    Green = 8'h85;    Blue = 8'h6b;
end 13'h104c:    begin Red = 8'h9c;    Green = 8'h8a;    Blue = 8'h69;
end 13'h104d:    begin Red = 8'ha0;    Green = 8'h8e;    Blue = 8'h69;
end 13'h104e:    begin Red = 8'hbc;    Green = 8'hb9;    Blue = 8'haf;
end 13'h104f:    begin Red = 8'he1;    Green = 8'hbe;    Blue = 8'ha3;
end 13'h1050:    begin Red = 8'hde;    Green = 8'hbb;    Blue = 8'h97;
end 13'h1051:    begin Red = 8'he3;    Green = 8'hba;    Blue = 8'h9a;
end 13'h1052:    begin Red = 8'hdd;    Green = 8'hb7;    Blue = 8'h97;
end 13'h1053:    begin Red = 8'h9e;    Green = 8'h88;    Blue = 8'h66;
end 13'h1054:    begin Red = 8'hd9;    Green = 8'hbd;    Blue = 8'h9d;
end 13'h1055:    begin Red = 8'hda;    Green = 8'hc1;    Blue = 8'h9a;
end 13'h1056:    begin Red = 8'hce;    Green = 8'hca;    Blue = 8'hb7;
end 13'h1057:    begin Red = 8'hc3;    Green = 8'hc8;    Blue = 8'ha0;
end 13'h1058:    begin Red = 8'h9c;    Green = 8'h97;    Blue = 8'h82;
end 13'h1059:    begin Red = 8'he6;    Green = 8'hdb;    Blue = 8'hc4;
end 13'h105a:    begin Red = 8'hb7;    Green = 8'hb7;    Blue = 8'ha1;
end 13'h105b:    begin Red = 8'hc6;    Green = 8'hc0;    Blue = 8'hb3;
end 13'h105c:    begin Red = 8'hd2;    Green = 8'he1;    Blue = 8'hb3;
end 13'h105d:    begin Red = 8'hd0;    Green = 8'hd8;    Blue = 8'haf;
end 13'h105e:    begin Red = 8'hac;    Green = 8'haa;    Blue = 8'h8e;
end 13'h105f:    begin Red = 8'ha9;    Green = 8'h85;    Blue = 8'h6c;
end 13'h1060:    begin Red = 8'he8;    Green = 8'hcc;    Blue = 8'hac;
end 13'h1061:    begin Red = 8'hb3;    Green = 8'h9a;    Blue = 8'h75;
end 13'h1062:    begin Red = 8'hbc;    Green = 8'hb4;    Blue = 8'hab;
end 13'h1063:    begin Red = 8'hc3;    Green = 8'ha1;    Blue = 8'h8d;
end 13'h1064:    begin Red = 8'h6c;    Green = 8'h6a;    Blue = 8'h56;
end 13'h1065:    begin Red = 8'hba;    Green = 8'ha0;    Blue = 8'h85;
end 13'h1066:    begin Red = 8'hd9;    Green = 8'hb8;    Blue = 8'h95;
end 13'h1067:    begin Red = 8'he6;    Green = 8'hd4;    Blue = 8'hb3;
end 13'h1068:    begin Red = 8'ha2;    Green = 8'hbf;    Blue = 8'ha7;
end 13'h1069:    begin Red = 8'hd5;    Green = 8'hc9;    Blue = 8'hb2;
end 13'h106a:    begin Red = 8'h9a;    Green = 8'ha0;    Blue = 8'h90;
end 13'h106b:    begin Red = 8'hec;    Green = 8'hb0;    Blue = 8'h7d;
end 13'h106c:    begin Red = 8'hc5;    Green = 8'h8e;    Blue = 8'h6f;
end 13'h106d:    begin Red = 8'hd3;    Green = 8'hd4;    Blue = 8'hbb;
end 13'h106e:    begin Red = 8'hc2;    Green = 8'h94;    Blue = 8'h74;
end 13'h106f:    begin Red = 8'hf9;    Green = 8'haf;    Blue = 8'h8c;
end 13'h1070:    begin Red = 8'hcd;    Green = 8'ha7;    Blue = 8'h83;
end 13'h1071:    begin Red = 8'haa;    Green = 8'h90;    Blue = 8'h67;
end 13'h1072:    begin Red = 8'hd5;    Green = 8'hc1;    Blue = 8'ha0;
end 13'h1073:    begin Red = 8'ha8;    Green = 8'h93;    Blue = 8'h6d;
end 13'h1074:    begin Red = 8'hd5;    Green = 8'hc0;    Blue = 8'ha4;
end 13'h1075:    begin Red = 8'hba;    Green = 8'hb2;    Blue = 8'ha8;
end 13'h1076:    begin Red = 8'hb7;    Green = 8'h9c;    Blue = 8'h80;
end 13'h1077:    begin Red = 8'ha9;    Green = 8'h94;    Blue = 8'h71;
end 13'h1078:    begin Red = 8'ha5;    Green = 8'hb4;    Blue = 8'ha3;
end 13'h1079:    begin Red = 8'hea;    Green = 8'hdc;    Blue = 8'hcf;
end 13'h107a:    begin Red = 8'he9;    Green = 8'he6;    Blue = 8'hca;
end 13'h107b:    begin Red = 8'hf7;    Green = 8'haf;    Blue = 8'h81;
end 13'h107c:    begin Red = 8'hf0;    Green = 8'hb1;    Blue = 8'h84;
end 13'h107d:    begin Red = 8'hce;    Green = 8'hdf;    Blue = 8'hc1;
end 13'h107e:    begin Red = 8'ha3;    Green = 8'haf;    Blue = 8'h88;
end 13'h107f:    begin Red = 8'hbf;    Green = 8'h98;    Blue = 8'h7f;
end 13'h1080:    begin Red = 8'hb4;    Green = 8'hc2;    Blue = 8'ha5;
end 13'h1081:    begin Red = 8'hb2;    Green = 8'h93;    Blue = 8'h78;
end 13'h1082:    begin Red = 8'he2;    Green = 8'hd0;    Blue = 8'hab;
end 13'h1083:    begin Red = 8'hd6;    Green = 8'hb7;    Blue = 8'h94;
end 13'h1084:    begin Red = 8'h65;    Green = 8'h60;    Blue = 8'h56;
end 13'h1085:    begin Red = 8'he1;    Green = 8'hd3;    Blue = 8'hc5;
end 13'h1086:    begin Red = 8'hde;    Green = 8'h9d;    Blue = 8'h71;
end 13'h1087:    begin Red = 8'hb8;    Green = 8'h9b;    Blue = 8'h77;
end 13'h1088:    begin Red = 8'hc9;    Green = 8'hcf;    Blue = 8'hb2;
end 13'h1089:    begin Red = 8'hb9;    Green = 8'h97;    Blue = 8'h7b;
end 13'h108a:    begin Red = 8'h95;    Green = 8'h7f;    Blue = 8'h61;
end 13'h108b:    begin Red = 8'ha7;    Green = 8'h90;    Blue = 8'h6e;
end 13'h108c:    begin Red = 8'hb9;    Green = 8'haf;    Blue = 8'ha7;
end 13'h108d:    begin Red = 8'h6e;    Green = 8'h62;    Blue = 8'h51;
end 13'h108e:    begin Red = 8'h62;    Green = 8'h54;    Blue = 8'h4c;
end 13'h108f:    begin Red = 8'h5f;    Green = 8'h50;    Blue = 8'h4b;
end 13'h1090:    begin Red = 8'h5d;    Green = 8'h4d;    Blue = 8'h4c;
end 13'h1091:    begin Red = 8'hd8;    Green = 8'hb8;    Blue = 8'h9b;
end 13'h1092:    begin Red = 8'hd0;    Green = 8'h84;    Blue = 8'h5e;
end 13'h1093:    begin Red = 8'he0;    Green = 8'hac;    Blue = 8'h8c;
end 13'h1094:    begin Red = 8'hc8;    Green = 8'hc5;    Blue = 8'hae;
end 13'h1095:    begin Red = 8'hc7;    Green = 8'h91;    Blue = 8'h3e;
end 13'h1096:    begin Red = 8'hd2;    Green = 8'h9a;    Blue = 8'h47;
end 13'h1097:    begin Red = 8'hcf;    Green = 8'h98;    Blue = 8'h46;
end 13'h1098:    begin Red = 8'hd5;    Green = 8'h99;    Blue = 8'h3e;
end 13'h1099:    begin Red = 8'hac;    Green = 8'h80;    Blue = 8'h5d;
end 13'h109a:    begin Red = 8'h77;    Green = 8'h9f;    Blue = 8'h75;
end 13'h109b:    begin Red = 8'h86;    Green = 8'hb7;    Blue = 8'h82;
end 13'h109c:    begin Red = 8'hdb;    Green = 8'he0;    Blue = 8'hc2;
end 13'h109d:    begin Red = 8'h7a;    Green = 8'h9f;    Blue = 8'h6c;
end 13'h109e:    begin Red = 8'h7f;    Green = 8'h96;    Blue = 8'h69;
end 13'h109f:    begin Red = 8'h84;    Green = 8'hb3;    Blue = 8'h7a;
end 13'h10a0:    begin Red = 8'hdc;    Green = 8'hc9;    Blue = 8'hac;
end 13'h10a1:    begin Red = 8'hd9;    Green = 8'hbb;    Blue = 8'h98;
end 13'h10a2:    begin Red = 8'hd2;    Green = 8'hbf;    Blue = 8'h96;
end 13'h10a3:    begin Red = 8'hcf;    Green = 8'hd2;    Blue = 8'hb9;
end 13'h10a4:    begin Red = 8'hd1;    Green = 8'hd4;    Blue = 8'hb8;
end 13'h10a5:    begin Red = 8'hc8;    Green = 8'h84;    Blue = 8'h5b;
end 13'h10a6:    begin Red = 8'heb;    Green = 8'had;    Blue = 8'h7c;
end 13'h10a7:    begin Red = 8'hf2;    Green = 8'ha7;    Blue = 8'h7e;
end 13'h10a8:    begin Red = 8'he4;    Green = 8'hb3;    Blue = 8'h78;
end 13'h10a9:    begin Red = 8'hec;    Green = 8'haf;    Blue = 8'h8c;
end 13'h10aa:    begin Red = 8'hf1;    Green = 8'hae;    Blue = 8'h83;
end 13'h10ab:    begin Red = 8'he1;    Green = 8'hea;    Blue = 8'hd7;
end 13'h10ac:    begin Red = 8'he2;    Green = 8'he6;    Blue = 8'hd0;
end 13'h10ad:    begin Red = 8'hd5;    Green = 8'hd4;    Blue = 8'hbe;
end 13'h10ae:    begin Red = 8'he7;    Green = 8'hb2;    Blue = 8'h88;
end 13'h10af:    begin Red = 8'hc5;    Green = 8'h9b;    Blue = 8'h76;
end 13'h10b0:    begin Red = 8'ha2;    Green = 8'haf;    Blue = 8'h99;
end 13'h10b1:    begin Red = 8'hc7;    Green = 8'h91;    Blue = 8'h70;
end 13'h10b2:    begin Red = 8'he5;    Green = 8'haf;    Blue = 8'h92;
end 13'h10b3:    begin Red = 8'hc9;    Green = 8'h94;    Blue = 8'h3a;
end 13'h10b4:    begin Red = 8'hca;    Green = 8'h9c;    Blue = 8'h42;
end 13'h10b5:    begin Red = 8'h8c;    Green = 8'hb7;    Blue = 8'h86;
end 13'h10b6:    begin Red = 8'ha6;    Green = 8'hab;    Blue = 8'h8e;
end 13'h10b7:    begin Red = 8'h79;    Green = 8'ha1;    Blue = 8'h71;
end 13'h10b8:    begin Red = 8'h8f;    Green = 8'hb6;    Blue = 8'h8a;
end 13'h10b9:    begin Red = 8'hcf;    Green = 8'hd3;    Blue = 8'hb3;
end 13'h10ba:    begin Red = 8'hcc;    Green = 8'hb9;    Blue = 8'h9b;
end 13'h10bb:    begin Red = 8'ha9;    Green = 8'h91;    Blue = 8'h73;
end 13'h10bc:    begin Red = 8'hcd;    Green = 8'hba;    Blue = 8'h9f;
end 13'h10bd:    begin Red = 8'hb5;    Green = 8'ha7;    Blue = 8'h88;
end 13'h10be:    begin Red = 8'h79;    Green = 8'h68;    Blue = 8'h55;
end 13'h10bf:    begin Red = 8'h73;    Green = 8'h61;    Blue = 8'h4f;
end 13'h10c0:    begin Red = 8'h6b;    Green = 8'h5d;    Blue = 8'h51;
end 13'h10c1:    begin Red = 8'h65;    Green = 8'h57;    Blue = 8'h51;
end 13'h10c2:    begin Red = 8'hcb;    Green = 8'hb0;    Blue = 8'h8c;
end 13'h10c3:    begin Red = 8'hc3;    Green = 8'hc2;    Blue = 8'hb6;
end 13'h10c4:    begin Red = 8'h86;    Green = 8'h84;    Blue = 8'h65;
end 13'h10c5:    begin Red = 8'h89;    Green = 8'h84;    Blue = 8'h71;
end 13'h10c6:    begin Red = 8'ha0;    Green = 8'h8b;    Blue = 8'h7c;
end 13'h10c7:    begin Red = 8'hc9;    Green = 8'h90;    Blue = 8'h5f;
end 13'h10c8:    begin Red = 8'he9;    Green = 8'hae;    Blue = 8'h8a;
end 13'h10c9:    begin Red = 8'he5;    Green = 8'hb3;    Blue = 8'h7c;
end 13'h10ca:    begin Red = 8'he2;    Green = 8'ha3;    Blue = 8'h75;
end 13'h10cb:    begin Red = 8'hea;    Green = 8'hdc;    Blue = 8'hc9;
end 13'h10cc:    begin Red = 8'h72;    Green = 8'h6d;    Blue = 8'h5a;
end 13'h10cd:    begin Red = 8'hc5;    Green = 8'hcb;    Blue = 8'ha4;
end 13'h10ce:    begin Red = 8'hec;    Green = 8'hac;    Blue = 8'h82;
end 13'h10cf:    begin Red = 8'hec;    Green = 8'ha6;    Blue = 8'h88;
end 13'h10d0:    begin Red = 8'he9;    Green = 8'hb3;    Blue = 8'h8c;
end 13'h10d1:    begin Red = 8'hf1;    Green = 8'hac;    Blue = 8'h4f;
end 13'h10d2:    begin Red = 8'hc7;    Green = 8'h93;    Blue = 8'h4b;
end 13'h10d3:    begin Red = 8'hce;    Green = 8'h98;    Blue = 8'h4b;
end 13'h10d4:    begin Red = 8'h9f;    Green = 8'h9c;    Blue = 8'h82;
end 13'h10d5:    begin Red = 8'hb5;    Green = 8'hab;    Blue = 8'ha3;
end 13'h10d6:    begin Red = 8'hc3;    Green = 8'ha2;    Blue = 8'h7c;
end 13'h10d7:    begin Red = 8'hb0;    Green = 8'h98;    Blue = 8'h7c;
end 13'h10d8:    begin Red = 8'h56;    Green = 8'h4f;    Blue = 8'h4b;
end 13'h10d9:    begin Red = 8'hcd;    Green = 8'haf;    Blue = 8'h90;
end 13'h10da:    begin Red = 8'hd2;    Green = 8'hbe;    Blue = 8'ha5;
end 13'h10db:    begin Red = 8'hc5;    Green = 8'hc7;    Blue = 8'ha7;
end 13'h10dc:    begin Red = 8'ha9;    Green = 8'h8e;    Blue = 8'h6a;
end 13'h10dd:    begin Red = 8'hc7;    Green = 8'hc7;    Blue = 8'hb1;
end 13'h10de:    begin Red = 8'hda;    Green = 8'hd5;    Blue = 8'hbe;
end 13'h10df:    begin Red = 8'hdd;    Green = 8'hf0;    Blue = 8'hf9;
end 13'h10e0:    begin Red = 8'hc0;    Green = 8'hc3;    Blue = 8'hae;
end 13'h10e1:    begin Red = 8'hc3;    Green = 8'hcb;    Blue = 8'hb2;
end 13'h10e2:    begin Red = 8'hc4;    Green = 8'hc7;    Blue = 8'haf;
end 13'h10e3:    begin Red = 8'hc1;    Green = 8'hc6;    Blue = 8'ha9;
end 13'h10e4:    begin Red = 8'h85;    Green = 8'h80;    Blue = 8'h6d;
end 13'h10e5:    begin Red = 8'hbd;    Green = 8'hc3;    Blue = 8'h9a;
end 13'h10e6:    begin Red = 8'ha2;    Green = 8'h96;    Blue = 8'h85;
end 13'h10e7:    begin Red = 8'hd5;    Green = 8'he7;    Blue = 8'hc4;
end 13'h10e8:    begin Red = 8'hac;    Green = 8'hac;    Blue = 8'h87;
end 13'h10e9:    begin Red = 8'ha5;    Green = 8'hb6;    Blue = 8'h95;
end 13'h10ea:    begin Red = 8'ha7;    Green = 8'h84;    Blue = 8'h69;
end 13'h10eb:    begin Red = 8'hf4;    Green = 8'haf;    Blue = 8'h42;
end 13'h10ec:    begin Red = 8'hd0;    Green = 8'h96;    Blue = 8'h4a;
end 13'h10ed:    begin Red = 8'hce;    Green = 8'hbd;    Blue = 8'ha0;
end 13'h10ee:    begin Red = 8'hfb;    Green = 8'he9;    Blue = 8'hc8;
end 13'h10ef:    begin Red = 8'h63;    Green = 8'h55;    Blue = 8'h4f;
end 13'h10f0:    begin Red = 8'h60;    Green = 8'h4b;    Blue = 8'h4e;
end 13'h10f1:    begin Red = 8'hae;    Green = 8'h99;    Blue = 8'h84;
end 13'h10f2:    begin Red = 8'ha5;    Green = 8'h95;    Blue = 8'h6d;
end 13'h10f3:    begin Red = 8'he0;    Green = 8'hd3;    Blue = 8'hc1;
end 13'h10f4:    begin Red = 8'hbf;    Green = 8'hd1;    Blue = 8'ha0;
end 13'h10f5:    begin Red = 8'hcf;    Green = 8'h98;    Blue = 8'h77;
end 13'h10f6:    begin Red = 8'hcd;    Green = 8'h99;    Blue = 8'h79;
end 13'h10f7:    begin Red = 8'hf2;    Green = 8'hb0;    Blue = 8'h47;
end 13'h10f8:    begin Red = 8'hb9;    Green = 8'hcb;    Blue = 8'haa;
end 13'h10f9:    begin Red = 8'h90;    Green = 8'h8b;    Blue = 8'h71;
end 13'h10fa:    begin Red = 8'hf1;    Green = 8'hd4;    Blue = 8'hac;
end 13'h10fb:    begin Red = 8'hd7;    Green = 8'hc0;    Blue = 8'h8c;
end 13'h10fc:    begin Red = 8'hd7;    Green = 8'hc1;    Blue = 8'h90;
end 13'h10fd:    begin Red = 8'hfb;    Green = 8'he0;    Blue = 8'hb1;
end 13'h10fe:    begin Red = 8'hd9;    Green = 8'hba;    Blue = 8'h8b;
end 13'h10ff:    begin Red = 8'hfa;    Green = 8'hde;    Blue = 8'hae;
end 13'h1100:    begin Red = 8'hcc;    Green = 8'hbd;    Blue = 8'h9d;
end 13'h1101:    begin Red = 8'hef;    Green = 8'hd9;    Blue = 8'haa;
end 13'h1102:    begin Red = 8'h83;    Green = 8'h6d;    Blue = 8'h56;
end 13'h1103:    begin Red = 8'h6c;    Green = 8'h5a;    Blue = 8'h4f;
end 13'h1104:    begin Red = 8'h47;    Green = 8'h38;    Blue = 8'h34;
end 13'h1105:    begin Red = 8'hee;    Green = 8'hd2;    Blue = 8'haa;
end 13'h1106:    begin Red = 8'hd9;    Green = 8'hb7;    Blue = 8'h87;
end 13'h1107:    begin Red = 8'hd5;    Green = 8'hb6;    Blue = 8'h87;
end 13'h1108:    begin Red = 8'hf0;    Green = 8'hd1;    Blue = 8'ha3;
end 13'h1109:    begin Red = 8'hd4;    Green = 8'hb8;    Blue = 8'h89;
end 13'h110a:    begin Red = 8'hfd;    Green = 8'hea;    Blue = 8'hbf;
end 13'h110b:    begin Red = 8'hfb;    Green = 8'he2;    Blue = 8'hbe;
end 13'h110c:    begin Red = 8'he8;    Green = 8'hd5;    Blue = 8'hb7;
end 13'h110d:    begin Red = 8'h87;    Green = 8'h72;    Blue = 8'h5d;
end 13'h110e:    begin Red = 8'hcb;    Green = 8'hb3;    Blue = 8'h87;
end 13'h110f:    begin Red = 8'hd4;    Green = 8'hbc;    Blue = 8'h8c;
end 13'h1110:    begin Red = 8'h3c;    Green = 8'h34;    Blue = 8'h27;
end 13'h1111:    begin Red = 8'h3e;    Green = 8'h37;    Blue = 8'h27;
end 13'h1112:    begin Red = 8'h3e;    Green = 8'h38;    Blue = 8'h20;
end 13'h1113:    begin Red = 8'hfa;    Green = 8'hcd;    Blue = 8'ha4;
end 13'h1114:    begin Red = 8'h9c;    Green = 8'h7c;    Blue = 8'h59;
end 13'h1115:    begin Red = 8'heb;    Green = 8'ha3;    Blue = 8'h72;
end 13'h1116:    begin Red = 8'he7;    Green = 8'he5;    Blue = 8'hcc;
end 13'h1117:    begin Red = 8'hf8;    Green = 8'hf9;    Blue = 8'he0;
end 13'h1118:    begin Red = 8'h80;    Green = 8'h80;    Blue = 8'h68;
end 13'h1119:    begin Red = 8'h85;    Green = 8'h84;    Blue = 8'h6c;
end 13'h111a:    begin Red = 8'hb8;    Green = 8'hbe;    Blue = 8'h96;
end 13'h111b:    begin Red = 8'heb;    Green = 8'h9f;    Blue = 8'h34;
end 13'h111c:    begin Red = 8'heb;    Green = 8'ha8;    Blue = 8'h4c;
end 13'h111d:    begin Red = 8'he3;    Green = 8'hac;    Blue = 8'h4f;
end 13'h111e:    begin Red = 8'he6;    Green = 8'hd3;    Blue = 8'ha9;
end 13'h111f:    begin Red = 8'hd8;    Green = 8'hbd;    Blue = 8'h90;
end 13'h1120:    begin Red = 8'hf5;    Green = 8'hd7;    Blue = 8'hb1;
end 13'h1121:    begin Red = 8'h81;    Green = 8'h71;    Blue = 8'h58;
end 13'h1122:    begin Red = 8'hc1;    Green = 8'hb2;    Blue = 8'h98;
end 13'h1123:    begin Red = 8'hac;    Green = 8'ha4;    Blue = 8'h9d;
end 13'h1124:    begin Red = 8'h4a;    Green = 8'h3f;    Blue = 8'h34;
end 13'h1125:    begin Red = 8'hf3;    Green = 8'hd2;    Blue = 8'haf;
end 13'h1126:    begin Red = 8'hd1;    Green = 8'hb7;    Blue = 8'h84;
end 13'h1127:    begin Red = 8'hdb;    Green = 8'hbf;    Blue = 8'h8f;
end 13'h1128:    begin Red = 8'hff;    Green = 8'hf4;    Blue = 8'hc6;
end 13'h1129:    begin Red = 8'hff;    Green = 8'hfd;    Blue = 8'hc9;
end 13'h112a:    begin Red = 8'hd7;    Green = 8'hd8;    Blue = 8'hb8;
end 13'h112b:    begin Red = 8'hfe;    Green = 8'hbb;    Blue = 8'h8c;
end 13'h112c:    begin Red = 8'hf7;    Green = 8'hbf;    Blue = 8'h90;
end 13'h112d:    begin Red = 8'hff;    Green = 8'hb6;    Blue = 8'h85;
end 13'h112e:    begin Red = 8'h98;    Green = 8'h90;    Blue = 8'h8c;
end 13'h112f:    begin Red = 8'h9a;    Green = 8'h91;    Blue = 8'h8e;
end 13'h1130:    begin Red = 8'h95;    Green = 8'h93;    Blue = 8'h8f;
end 13'h1131:    begin Red = 8'h88;    Green = 8'h6d;    Blue = 8'h4a;
end 13'h1132:    begin Red = 8'h94;    Green = 8'h8a;    Blue = 8'h6c;
end 13'h1133:    begin Red = 8'hd5;    Green = 8'h8d;    Blue = 8'h5d;
end 13'h1134:    begin Red = 8'hff;    Green = 8'hbe;    Blue = 8'h89;
end 13'h1135:    begin Red = 8'hff;    Green = 8'hc0;    Blue = 8'h8c;
end 13'h1136:    begin Red = 8'hff;    Green = 8'hbd;    Blue = 8'h84;
end 13'h1137:    begin Red = 8'he2;    Green = 8'he5;    Blue = 8'hd9;
end 13'h1138:    begin Red = 8'hd6;    Green = 8'hcb;    Blue = 8'hb0;
end 13'h1139:    begin Red = 8'hee;    Green = 8'ha1;    Blue = 8'h37;
end 13'h113a:    begin Red = 8'hfd;    Green = 8'hb2;    Blue = 8'h4e;
end 13'h113b:    begin Red = 8'hf5;    Green = 8'hb3;    Blue = 8'h4a;
end 13'h113c:    begin Red = 8'hd2;    Green = 8'h97;    Blue = 8'h40;
end 13'h113d:    begin Red = 8'hac;    Green = 8'h8c;    Blue = 8'h5d;
end 13'h113e:    begin Red = 8'h63;    Green = 8'h68;    Blue = 8'h60;
end 13'h113f:    begin Red = 8'hcf;    Green = 8'hb3;    Blue = 8'h83;
end 13'h1140:    begin Red = 8'he2;    Green = 8'hd2;    Blue = 8'haf;
end 13'h1141:    begin Red = 8'h8e;    Green = 8'h7f;    Blue = 8'h67;
end 13'h1142:    begin Red = 8'hf2;    Green = 8'hd7;    Blue = 8'haa;
end 13'h1143:    begin Red = 8'hea;    Green = 8'hcf;    Blue = 8'ha0;
end 13'h1144:    begin Red = 8'hfb;    Green = 8'hdc;    Blue = 8'ha5;
end 13'h1145:    begin Red = 8'hed;    Green = 8'hae;    Blue = 8'h87;
end 13'h1146:    begin Red = 8'h90;    Green = 8'h80;    Blue = 8'h81;
end 13'h1147:    begin Red = 8'h9a;    Green = 8'h90;    Blue = 8'h83;
end 13'h1148:    begin Red = 8'h9c;    Green = 8'h92;    Blue = 8'h85;
end 13'h1149:    begin Red = 8'hcf;    Green = 8'h8c;    Blue = 8'h58;
end 13'h114a:    begin Red = 8'heb;    Green = 8'hdc;    Blue = 8'hc3;
end 13'h114b:    begin Red = 8'hca;    Green = 8'hc2;    Blue = 8'haa;
end 13'h114c:    begin Red = 8'hc4;    Green = 8'hbb;    Blue = 8'haa;
end 13'h114d:    begin Red = 8'hed;    Green = 8'hae;    Blue = 8'h4f;
end 13'h114e:    begin Red = 8'hfd;    Green = 8'hb3;    Blue = 8'h42;
end 13'h114f:    begin Red = 8'hfb;    Green = 8'hb5;    Blue = 8'h4b;
end 13'h1150:    begin Red = 8'hdc;    Green = 8'h9b;    Blue = 8'h45;
end 13'h1151:    begin Red = 8'h75;    Green = 8'h7e;    Blue = 8'h65;
end 13'h1152:    begin Red = 8'h66;    Green = 8'h74;    Blue = 8'h59;
end 13'h1153:    begin Red = 8'h65;    Green = 8'h74;    Blue = 8'h64;
end 13'h1154:    begin Red = 8'h71;    Green = 8'h7f;    Blue = 8'h64;
end 13'h1155:    begin Red = 8'had;    Green = 8'ha0;    Blue = 8'ha0;
end 13'h1156:    begin Red = 8'ha0;    Green = 8'h8d;    Blue = 8'h7f;
end 13'h1157:    begin Red = 8'hc5;    Green = 8'haa;    Blue = 8'h85;
end 13'h1158:    begin Red = 8'ha3;    Green = 8'hac;    Blue = 8'h90;
end 13'h1159:    begin Red = 8'hd9;    Green = 8'hc8;    Blue = 8'hab;
end 13'h115a:    begin Red = 8'hb8;    Green = 8'hb8;    Blue = 8'h9c;
end 13'h115b:    begin Red = 8'h8e;    Green = 8'h84;    Blue = 8'h7d;
end 13'h115c:    begin Red = 8'hcb;    Green = 8'hae;    Blue = 8'h76;
end 13'h115d:    begin Red = 8'hc7;    Green = 8'hac;    Blue = 8'h71;
end 13'h115e:    begin Red = 8'hca;    Green = 8'ha8;    Blue = 8'h6c;
end 13'h115f:    begin Red = 8'hc9;    Green = 8'hac;    Blue = 8'h6e;
end 13'h1160:    begin Red = 8'hc7;    Green = 8'h86;    Blue = 8'h64;
end 13'h1161:    begin Red = 8'hee;    Green = 8'hac;    Blue = 8'h78;
end 13'h1162:    begin Red = 8'hd5;    Green = 8'h9b;    Blue = 8'h74;
end 13'h1163:    begin Red = 8'he5;    Green = 8'had;    Blue = 8'h8c;
end 13'h1164:    begin Red = 8'heb;    Green = 8'hd6;    Blue = 8'hcc;
end 13'h1165:    begin Red = 8'hc0;    Green = 8'h9b;    Blue = 8'h75;
end 13'h1166:    begin Red = 8'hd1;    Green = 8'he3;    Blue = 8'hc2;
end 13'h1167:    begin Red = 8'hbe;    Green = 8'h98;    Blue = 8'h74;
end 13'h1168:    begin Red = 8'h67;    Green = 8'h56;    Blue = 8'h3e;
end 13'h1169:    begin Red = 8'h75;    Green = 8'h65;    Blue = 8'h58;
end 13'h116a:    begin Red = 8'hd8;    Green = 8'hc5;    Blue = 8'ha8;
end 13'h116b:    begin Red = 8'h9e;    Green = 8'h96;    Blue = 8'h95;
end 13'h116c:    begin Red = 8'h5a;    Green = 8'h4d;    Blue = 8'h3a;
end 13'h116d:    begin Red = 8'h53;    Green = 8'h46;    Blue = 8'h3a;
end 13'h116e:    begin Red = 8'h45;    Green = 8'h34;    Blue = 8'h34;
end 13'h116f:    begin Red = 8'hd5;    Green = 8'hc3;    Blue = 8'ha9;
end 13'h1170:    begin Red = 8'h51;    Green = 8'h4d;    Blue = 8'h34;
end 13'h1171:    begin Red = 8'ha4;    Green = 8'h9a;    Blue = 8'h95;
end 13'h1172:    begin Red = 8'hf9;    Green = 8'hff;    Blue = 8'hf9;
end 13'h1173:    begin Red = 8'hfb;    Green = 8'hfc;    Blue = 8'hed;
end 13'h1174:    begin Red = 8'hc9;    Green = 8'ha7;    Blue = 8'h58;
end 13'h1175:    begin Red = 8'hc3;    Green = 8'haa;    Blue = 8'h68;
end 13'h1176:    begin Red = 8'hcf;    Green = 8'hb2;    Blue = 8'h6c;
end 13'h1177:    begin Red = 8'hcb;    Green = 8'haf;    Blue = 8'h6c;
end 13'h1178:    begin Red = 8'hd1;    Green = 8'hb5;    Blue = 8'h74;
end 13'h1179:    begin Red = 8'hf1;    Green = 8'ha7;    Blue = 8'h77;
end 13'h117a:    begin Red = 8'hee;    Green = 8'ha8;    Blue = 8'h82;
end 13'h117b:    begin Red = 8'hf7;    Green = 8'ha9;    Blue = 8'h78;
end 13'h117c:    begin Red = 8'hcb;    Green = 8'h90;    Blue = 8'h6b;
end 13'h117d:    begin Red = 8'hdc;    Green = 8'hed;    Blue = 8'hd4;
end 13'h117e:    begin Red = 8'hdf;    Green = 8'heb;    Blue = 8'hdc;
end 13'h117f:    begin Red = 8'h89;    Green = 8'h8f;    Blue = 8'h75;
end 13'h1180:    begin Red = 8'he7;    Green = 8'hc7;    Blue = 8'h96;
end 13'h1181:    begin Red = 8'hea;    Green = 8'hca;    Blue = 8'h99;
end 13'h1182:    begin Red = 8'he6;    Green = 8'hc7;    Blue = 8'h9b;
end 13'h1183:    begin Red = 8'hea;    Green = 8'hcb;    Blue = 8'h95;
end 13'h1184:    begin Red = 8'hc9;    Green = 8'ha7;    Blue = 8'h7a;
end 13'h1185:    begin Red = 8'hc9;    Green = 8'haa;    Blue = 8'h7e;
end 13'h1186:    begin Red = 8'hc6;    Green = 8'ha4;    Blue = 8'h77;
end 13'h1187:    begin Red = 8'he8;    Green = 8'hc9;    Blue = 8'h90;
end 13'h1188:    begin Red = 8'hea;    Green = 8'hc2;    Blue = 8'h9f;
end 13'h1189:    begin Red = 8'hdb;    Green = 8'hcb;    Blue = 8'h97;
end 13'h118a:    begin Red = 8'he4;    Green = 8'hc9;    Blue = 8'h9c;
end 13'h118b:    begin Red = 8'he4;    Green = 8'hc5;    Blue = 8'h99;
end 13'h118c:    begin Red = 8'he6;    Green = 8'hc8;    Blue = 8'h92;
end 13'h118d:    begin Red = 8'he6;    Green = 8'hc2;    Blue = 8'h8e;
end 13'h118e:    begin Red = 8'hcc;    Green = 8'hac;    Blue = 8'h86;
end 13'h118f:    begin Red = 8'hff;    Green = 8'hd4;    Blue = 8'h9f;
end 13'h1190:    begin Red = 8'hec;    Green = 8'hcd;    Blue = 8'h97;
end 13'h1191:    begin Red = 8'he4;    Green = 8'hc6;    Blue = 8'ha0;
end 13'h1192:    begin Red = 8'he7;    Green = 8'hc5;    Blue = 8'h9f;
end 13'h1193:    begin Red = 8'hde;    Green = 8'hc2;    Blue = 8'h90;
end 13'h1194:    begin Red = 8'he5;    Green = 8'hb0;    Blue = 8'h82;
end 13'h1195:    begin Red = 8'h90;    Green = 8'h86;    Blue = 8'h7b;
end 13'h1196:    begin Red = 8'hf9;    Green = 8'hea;    Blue = 8'hd2;
end 13'h1197:    begin Red = 8'hb1;    Green = 8'h9a;    Blue = 8'h65;
end 13'h1198:    begin Red = 8'hce;    Green = 8'hb1;    Blue = 8'h73;
end 13'h1199:    begin Red = 8'hcd;    Green = 8'hb3;    Blue = 8'h70;
end 13'h119a:    begin Red = 8'hac;    Green = 8'h94;    Blue = 8'h61;
end 13'h119b:    begin Red = 8'hbe;    Green = 8'hc9;    Blue = 8'hb4;
end 13'h119c:    begin Red = 8'hea;    Green = 8'ha5;    Blue = 8'h6e;
end 13'h119d:    begin Red = 8'hbf;    Green = 8'hc6;    Blue = 8'h9d;
end 13'h119e:    begin Red = 8'hc4;    Green = 8'hcb;    Blue = 8'ha9;
end 13'h119f:    begin Red = 8'hae;    Green = 8'h90;    Blue = 8'h6f;
end 13'h11a0:    begin Red = 8'h95;    Green = 8'h93;    Blue = 8'h77;
end 13'h11a1:    begin Red = 8'hcb;    Green = 8'haf;    Blue = 8'h7f;
end 13'h11a2:    begin Red = 8'hb3;    Green = 8'h92;    Blue = 8'h5c;
end 13'h11a3:    begin Red = 8'hb9;    Green = 8'h98;    Blue = 8'h63;
end 13'h11a4:    begin Red = 8'hd3;    Green = 8'hb2;    Blue = 8'h85;
end 13'h11a5:    begin Red = 8'h86;    Green = 8'h76;    Blue = 8'h5c;
end 13'h11a6:    begin Red = 8'h3b;    Green = 8'h2d;    Blue = 8'h2c;
end 13'h11a7:    begin Red = 8'h3b;    Green = 8'h29;    Blue = 8'h11;
end 13'h11a8:    begin Red = 8'h03;    Green = 8'h12;    Blue = 8'h68;
end 13'h11a9:    begin Red = 8'h42;    Green = 8'h39;    Blue = 8'h30;
end 13'h11aa:    begin Red = 8'h53;    Green = 8'h3b;    Blue = 8'h21;
end 13'h11ab:    begin Red = 8'h52;    Green = 8'h3b;    Blue = 8'h1b;
end 13'h11ac:    begin Red = 8'h3e;    Green = 8'h37;    Blue = 8'h2d;
end 13'h11ad:    begin Red = 8'h51;    Green = 8'h3d;    Blue = 8'h24;
end 13'h11ae:    begin Red = 8'h4c;    Green = 8'h3b;    Blue = 8'h1d;
end 13'h11af:    begin Red = 8'h40;    Green = 8'h34;    Blue = 8'h24;
end 13'h11b0:    begin Red = 8'h40;    Green = 8'h33;    Blue = 8'h20;
end 13'h11b1:    begin Red = 8'h40;    Green = 8'h3a;    Blue = 8'h2c;
end 13'h11b2:    begin Red = 8'h41;    Green = 8'h38;    Blue = 8'h29;
end 13'h11b3:    begin Red = 8'h40;    Green = 8'h32;    Blue = 8'h27;
end 13'h11b4:    begin Red = 8'hd1;    Green = 8'haf;    Blue = 8'h81;
end 13'h11b5:    begin Red = 8'hb7;    Green = 8'h95;    Blue = 8'h65;
end 13'h11b6:    begin Red = 8'hd2;    Green = 8'hb1;    Blue = 8'h88;
end 13'h11b7:    begin Red = 8'hb6;    Green = 8'h92;    Blue = 8'h62;
end 13'h11b8:    begin Red = 8'hcd;    Green = 8'hb5;    Blue = 8'h85;
end 13'h11b9:    begin Red = 8'h3b;    Green = 8'h32;    Blue = 8'h2b;
end 13'h11ba:    begin Red = 8'h2d;    Green = 8'h24;    Blue = 8'h1b;
end 13'h11bb:    begin Red = 8'h46;    Green = 8'h3d;    Blue = 8'h2e;
end 13'h11bc:    begin Red = 8'h89;    Green = 8'h66;    Blue = 8'h3c;
end 13'h11bd:    begin Red = 8'h31;    Green = 8'h35;    Blue = 8'h34;
end 13'h11be:    begin Red = 8'h45;    Green = 8'h38;    Blue = 8'h2f;
end 13'h11bf:    begin Red = 8'h61;    Green = 8'h4f;    Blue = 8'h37;
end 13'h11c0:    begin Red = 8'h67;    Green = 8'h4d;    Blue = 8'h3e;
end 13'h11c1:    begin Red = 8'h5b;    Green = 8'h3d;    Blue = 8'h19;
end 13'h11c2:    begin Red = 8'h47;    Green = 8'h33;    Blue = 8'h3e;
end 13'h11c3:    begin Red = 8'h04;    Green = 8'h72;    Blue = 8'hfd;
end 13'h11c4:    begin Red = 8'h41;    Green = 8'h39;    Blue = 8'h36;
end 13'h11c5:    begin Red = 8'h03;    Green = 8'h21;    Blue = 8'hdc;
end 13'h11c6:    begin Red = 8'h00;    Green = 8'h1b;    Blue = 8'h70;
end 13'h11c7:    begin Red = 8'hce;    Green = 8'hb1;    Blue = 8'h87;
end 13'h11c8:    begin Red = 8'hbb;    Green = 8'h95;    Blue = 8'h64;
end 13'h11c9:    begin Red = 8'hec;    Green = 8'hbf;    Blue = 8'h88;
end 13'h11ca:    begin Red = 8'h37;    Green = 8'h27;    Blue = 8'h2a;
end 13'h11cb:    begin Red = 8'h34;    Green = 8'h30;    Blue = 8'h25;
end 13'h11cc:    begin Red = 8'hda;    Green = 8'hda;    Blue = 8'hbc;
end 13'h11cd:    begin Red = 8'hbf;    Green = 8'h9b;    Blue = 8'h8b;
end 13'h11ce:    begin Red = 8'h40;    Green = 8'h35;    Blue = 8'h31;
end 13'h11cf:    begin Red = 8'h59;    Green = 8'h4b;    Blue = 8'h31;
end 13'h11d0:    begin Red = 8'h55;    Green = 8'h44;    Blue = 8'h30;
end 13'h11d1:    begin Red = 8'h42;    Green = 8'h37;    Blue = 8'h33;
end 13'h11d2:    begin Red = 8'h50;    Green = 8'h44;    Blue = 8'h2e;
end 13'h11d3:    begin Red = 8'h30;    Green = 8'h2a;    Blue = 8'h2c;
end 13'h11d4:    begin Red = 8'h34;    Green = 8'h2d;    Blue = 8'h1d;
end 13'h11d5:    begin Red = 8'h5e;    Green = 8'h51;    Blue = 8'h40;
end 13'h11d6:    begin Red = 8'h43;    Green = 8'h36;    Blue = 8'h2d;
end 13'h11d7:    begin Red = 8'h3d;    Green = 8'h34;    Blue = 8'h2f;
end 13'h11d8:    begin Red = 8'h45;    Green = 8'h36;    Blue = 8'h17;
end 13'h11d9:    begin Red = 8'h45;    Green = 8'h3b;    Blue = 8'h31;
end 13'h11da:    begin Red = 8'h3d;    Green = 8'h39;    Blue = 8'h30;
end 13'h11db:    begin Red = 8'h03;    Green = 8'h52;    Blue = 8'hac;
end 13'h11dc:    begin Red = 8'h79;    Green = 8'h5f;    Blue = 8'h52;
end 13'h11dd:    begin Red = 8'h56;    Green = 8'h4f;    Blue = 8'h35;
end 13'h11de:    begin Red = 8'h52;    Green = 8'h4b;    Blue = 8'h2e;
end 13'h11df:    begin Red = 8'h55;    Green = 8'h42;    Blue = 8'h33;
end 13'h11e0:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'h99;
end 13'h11e1:    begin Red = 8'h02;    Green = 8'h91;    Blue = 8'h79;
end 13'h11e2:    begin Red = 8'hd5;    Green = 8'haf;    Blue = 8'h8b;
end 13'h11e3:    begin Red = 8'hc6;    Green = 8'hb9;    Blue = 8'h85;
end 13'h11e4:    begin Red = 8'hea;    Green = 8'hf9;    Blue = 8'he2;
end 13'h11e5:    begin Red = 8'hf1;    Green = 8'hf3;    Blue = 8'he2;
end 13'h11e6:    begin Red = 8'hef;    Green = 8'hf5;    Blue = 8'hda;
end 13'h11e7:    begin Red = 8'hf1;    Green = 8'hf6;    Blue = 8'hec;
end 13'h11e8:    begin Red = 8'h8c;    Green = 8'h6f;    Blue = 8'h43;
end 13'h11e9:    begin Red = 8'hf9;    Green = 8'hf0;    Blue = 8'hd6;
end 13'h11ea:    begin Red = 8'hd0;    Green = 8'hcf;    Blue = 8'hbf;
end 13'h11eb:    begin Red = 8'hcc;    Green = 8'hac;    Blue = 8'h6a;
end 13'h11ec:    begin Red = 8'hc8;    Green = 8'had;    Blue = 8'h75;
end 13'h11ed:    begin Red = 8'h83;    Green = 8'h7d;    Blue = 8'h7b;
end 13'h11ee:    begin Red = 8'haf;    Green = 8'h72;    Blue = 8'h5a;
end 13'h11ef:    begin Red = 8'ha7;    Green = 8'h74;    Blue = 8'h5a;
end 13'h11f0:    begin Red = 8'ha9;    Green = 8'h7a;    Blue = 8'h5a;
end 13'h11f1:    begin Red = 8'ha7;    Green = 8'h7a;    Blue = 8'h56;
end 13'h11f2:    begin Red = 8'ha7;    Green = 8'h76;    Blue = 8'h57;
end 13'h11f3:    begin Red = 8'h5a;    Green = 8'h4a;    Blue = 8'h3c;
end 13'h11f4:    begin Red = 8'h42;    Green = 8'h41;    Blue = 8'h34;
end 13'h11f5:    begin Red = 8'hc1;    Green = 8'h90;    Blue = 8'h6d;
end 13'h11f6:    begin Red = 8'hc2;    Green = 8'h88;    Blue = 8'h67;
end 13'h11f7:    begin Red = 8'h88;    Green = 8'h8c;    Blue = 8'h6e;
end 13'h11f8:    begin Red = 8'h7e;    Green = 8'h70;    Blue = 8'h66;
end 13'h11f9:    begin Red = 8'hfc;    Green = 8'hf7;    Blue = 8'hde;
end 13'h11fa:    begin Red = 8'hfe;    Green = 8'hf9;    Blue = 8'he0;
end 13'h11fb:    begin Red = 8'h9e;    Green = 8'h7f;    Blue = 8'h5d;
end 13'h11fc:    begin Red = 8'hbd;    Green = 8'h9f;    Blue = 8'h69;
end 13'h11fd:    begin Red = 8'h55;    Green = 8'h43;    Blue = 8'h39;
end 13'h11fe:    begin Red = 8'h5b;    Green = 8'h46;    Blue = 8'h27;
end 13'h11ff:    begin Red = 8'h53;    Green = 8'h49;    Blue = 8'h26;
end 13'h1200:    begin Red = 8'h6c;    Green = 8'h55;    Blue = 8'h33;
end 13'h1201:    begin Red = 8'h69;    Green = 8'h57;    Blue = 8'h31;
end 13'h1202:    begin Red = 8'h6d;    Green = 8'h5d;    Blue = 8'h39;
end 13'h1203:    begin Red = 8'h61;    Green = 8'h52;    Blue = 8'h33;
end 13'h1204:    begin Red = 8'h5b;    Green = 8'h4c;    Blue = 8'h2d;
end 13'h1205:    begin Red = 8'h56;    Green = 8'h4a;    Blue = 8'h3e;
end 13'h1206:    begin Red = 8'hc9;    Green = 8'hbb;    Blue = 8'h98;
end 13'h1207:    begin Red = 8'h3c;    Green = 8'h39;    Blue = 8'h28;
end 13'h1208:    begin Red = 8'h32;    Green = 8'h2b;    Blue = 8'h19;
end 13'h1209:    begin Red = 8'hb6;    Green = 8'ha8;    Blue = 8'h81;
end 13'h120a:    begin Red = 8'h65;    Green = 8'h54;    Blue = 8'h44;
end 13'h120b:    begin Red = 8'ha7;    Green = 8'h7d;    Blue = 8'h53;
end 13'h120c:    begin Red = 8'h4d;    Green = 8'h4a;    Blue = 8'h45;
end 13'h120d:    begin Red = 8'h5c;    Green = 8'h4b;    Blue = 8'h41;
end 13'h120e:    begin Red = 8'h7a;    Green = 8'h67;    Blue = 8'h46;
end 13'h120f:    begin Red = 8'h74;    Green = 8'h56;    Blue = 8'h20;
end 13'h1210:    begin Red = 8'h63;    Green = 8'h47;    Blue = 8'h22;
end 13'h1211:    begin Red = 8'h54;    Green = 8'h39;    Blue = 8'h24;
end 13'h1212:    begin Red = 8'h03;    Green = 8'h31;    Blue = 8'hc0;
end 13'h1213:    begin Red = 8'hc4;    Green = 8'ha0;    Blue = 8'h70;
end 13'h1214:    begin Red = 8'hd0;    Green = 8'hb4;    Blue = 8'h8d;
end 13'h1215:    begin Red = 8'hd6;    Green = 8'hb4;    Blue = 8'h8e;
end 13'h1216:    begin Red = 8'hed;    Green = 8'hc8;    Blue = 8'h94;
end 13'h1217:    begin Red = 8'h38;    Green = 8'h39;    Blue = 8'h34;
end 13'h1218:    begin Red = 8'hd9;    Green = 8'hdc;    Blue = 8'hb8;
end 13'h1219:    begin Red = 8'hcd;    Green = 8'hba;    Blue = 8'h8f;
end 13'h121a:    begin Red = 8'h6c;    Green = 8'h5b;    Blue = 8'h3d;
end 13'h121b:    begin Red = 8'h5e;    Green = 8'h52;    Blue = 8'h46;
end 13'h121c:    begin Red = 8'h6d;    Green = 8'h60;    Blue = 8'h3d;
end 13'h121d:    begin Red = 8'h49;    Green = 8'h41;    Blue = 8'h36;
end 13'h121e:    begin Red = 8'h40;    Green = 8'h30;    Blue = 8'h30;
end 13'h121f:    begin Red = 8'h4e;    Green = 8'h41;    Blue = 8'h38;
end 13'h1220:    begin Red = 8'h67;    Green = 8'h57;    Blue = 8'h4a;
end 13'h1221:    begin Red = 8'ha7;    Green = 8'h8d;    Blue = 8'h7c;
end 13'h1222:    begin Red = 8'h66;    Green = 8'h4d;    Blue = 8'h2e;
end 13'h1223:    begin Red = 8'h64;    Green = 8'h56;    Blue = 8'h49;
end 13'h1224:    begin Red = 8'h73;    Green = 8'h56;    Blue = 8'h36;
end 13'h1225:    begin Red = 8'h5d;    Green = 8'h51;    Blue = 8'h53;
end 13'h1226:    begin Red = 8'h57;    Green = 8'h49;    Blue = 8'h2f;
end 13'h1227:    begin Red = 8'h91;    Green = 8'h77;    Blue = 8'h52;
end 13'h1228:    begin Red = 8'hcf;    Green = 8'hb9;    Blue = 8'h8a;
end 13'h1229:    begin Red = 8'h47;    Green = 8'h37;    Blue = 8'h20;
end 13'h122a:    begin Red = 8'hd3;    Green = 8'hb2;    Blue = 8'h7d;
end 13'h122b:    begin Red = 8'h9f;    Green = 8'h90;    Blue = 8'h84;
end 13'h122c:    begin Red = 8'ha3;    Green = 8'h95;    Blue = 8'h6a;
end 13'h122d:    begin Red = 8'hca;    Green = 8'hac;    Blue = 8'h5b;
end 13'h122e:    begin Red = 8'hd2;    Green = 8'hb8;    Blue = 8'h76;
end 13'h122f:    begin Red = 8'ha4;    Green = 8'h8a;    Blue = 8'h53;
end 13'h1230:    begin Red = 8'haa;    Green = 8'h8d;    Blue = 8'h52;
end 13'h1231:    begin Red = 8'hd5;    Green = 8'hb5;    Blue = 8'h71;
end 13'h1232:    begin Red = 8'hd9;    Green = 8'hbc;    Blue = 8'h7d;
end 13'h1233:    begin Red = 8'hac;    Green = 8'h6c;    Blue = 8'h54;
end 13'h1234:    begin Red = 8'ha0;    Green = 8'h72;    Blue = 8'h46;
end 13'h1235:    begin Red = 8'hb6;    Green = 8'h7d;    Blue = 8'h59;
end 13'h1236:    begin Red = 8'hb7;    Green = 8'h7d;    Blue = 8'h55;
end 13'h1237:    begin Red = 8'he2;    Green = 8'ha4;    Blue = 8'h80;
end 13'h1238:    begin Red = 8'h87;    Green = 8'h7f;    Blue = 8'h69;
end 13'h1239:    begin Red = 8'hc2;    Green = 8'h8a;    Blue = 8'h5b;
end 13'h123a:    begin Red = 8'hc8;    Green = 8'h8e;    Blue = 8'h6a;
end 13'h123b:    begin Red = 8'hd9;    Green = 8'h9f;    Blue = 8'h76;
end 13'h123c:    begin Red = 8'hcc;    Green = 8'h98;    Blue = 8'h6d;
end 13'h123d:    begin Red = 8'hce;    Green = 8'h93;    Blue = 8'h61;
end 13'h123e:    begin Red = 8'hae;    Green = 8'h9e;    Blue = 8'h8b;
end 13'h123f:    begin Red = 8'hc8;    Green = 8'hcf;    Blue = 8'had;
end 13'h1240:    begin Red = 8'hde;    Green = 8'he5;    Blue = 8'hbf;
end 13'h1241:    begin Red = 8'ha7;    Green = 8'h80;    Blue = 8'h62;
end 13'h1242:    begin Red = 8'hdd;    Green = 8'hbc;    Blue = 8'h8f;
end 13'h1243:    begin Red = 8'hdc;    Green = 8'hbe;    Blue = 8'h8c;
end 13'h1244:    begin Red = 8'h4f;    Green = 8'h42;    Blue = 8'h22;
end 13'h1245:    begin Red = 8'h62;    Green = 8'h56;    Blue = 8'h3c;
end 13'h1246:    begin Red = 8'h53;    Green = 8'h44;    Blue = 8'h25;
end 13'h1247:    begin Red = 8'h6a;    Green = 8'h56;    Blue = 8'h35;
end 13'h1248:    begin Red = 8'h69;    Green = 8'h51;    Blue = 8'h2d;
end 13'h1249:    begin Red = 8'h5c;    Green = 8'h4d;    Blue = 8'h30;
end 13'h124a:    begin Red = 8'h30;    Green = 8'h27;    Blue = 8'h16;
end 13'h124b:    begin Red = 8'h59;    Green = 8'h49;    Blue = 8'h39;
end 13'h124c:    begin Red = 8'ha5;    Green = 8'h96;    Blue = 8'h75;
end 13'h124d:    begin Red = 8'h64;    Green = 8'h52;    Blue = 8'h3c;
end 13'h124e:    begin Red = 8'h64;    Green = 8'h51;    Blue = 8'h4a;
end 13'h124f:    begin Red = 8'h8c;    Green = 8'h6d;    Blue = 8'h51;
end 13'h1250:    begin Red = 8'h85;    Green = 8'h6c;    Blue = 8'h4e;
end 13'h1251:    begin Red = 8'h73;    Green = 8'h59;    Blue = 8'h26;
end 13'h1252:    begin Red = 8'h5d;    Green = 8'h41;    Blue = 8'h2c;
end 13'h1253:    begin Red = 8'h61;    Green = 8'h44;    Blue = 8'h26;
end 13'h1254:    begin Red = 8'h5c;    Green = 8'h42;    Blue = 8'h29;
end 13'h1255:    begin Red = 8'h03;    Green = 8'h41;    Blue = 8'hf0;
end 13'h1256:    begin Red = 8'ha4;    Green = 8'h81;    Blue = 8'h61;
end 13'h1257:    begin Red = 8'h5a;    Green = 8'h46;    Blue = 8'h3b;
end 13'h1258:    begin Red = 8'h62;    Green = 8'h53;    Blue = 8'h3e;
end 13'h1259:    begin Red = 8'h55;    Green = 8'h48;    Blue = 8'h28;
end 13'h125a:    begin Red = 8'h64;    Green = 8'h55;    Blue = 8'h36;
end 13'h125b:    begin Red = 8'h5c;    Green = 8'h48;    Blue = 8'h2d;
end 13'h125c:    begin Red = 8'h62;    Green = 8'h51;    Blue = 8'h47;
end 13'h125d:    begin Red = 8'h57;    Green = 8'h49;    Blue = 8'h22;
end 13'h125e:    begin Red = 8'h66;    Green = 8'h52;    Blue = 8'h47;
end 13'h125f:    begin Red = 8'h42;    Green = 8'h37;    Blue = 8'h23;
end 13'h1260:    begin Red = 8'h47;    Green = 8'h34;    Blue = 8'h23;
end 13'h1261:    begin Red = 8'h96;    Green = 8'h7e;    Blue = 8'h56;
end 13'h1262:    begin Red = 8'hf1;    Green = 8'he7;    Blue = 8'hd8;
end 13'h1263:    begin Red = 8'h8f;    Green = 8'h7d;    Blue = 8'h53;
end 13'h1264:    begin Red = 8'h9d;    Green = 8'h87;    Blue = 8'h5f;
end 13'h1265:    begin Red = 8'hdb;    Green = 8'hd4;    Blue = 8'hc8;
end 13'h1266:    begin Red = 8'h82;    Green = 8'h73;    Blue = 8'h6d;
end 13'h1267:    begin Red = 8'h85;    Green = 8'h84;    Blue = 8'h75;
end 13'h1268:    begin Red = 8'h50;    Green = 8'h3d;    Blue = 8'h34;
end 13'h1269:    begin Red = 8'h83;    Green = 8'h7f;    Blue = 8'h65;
end 13'h126a:    begin Red = 8'hf6;    Green = 8'hf1;    Blue = 8'hdc;
end 13'h126b:    begin Red = 8'hd3;    Green = 8'hb0;    Blue = 8'h93;
end 13'h126c:    begin Red = 8'hb0;    Green = 8'hb1;    Blue = 8'h96;
end 13'h126d:    begin Red = 8'h53;    Green = 8'h43;    Blue = 8'h2a;
end 13'h126e:    begin Red = 8'h5d;    Green = 8'h50;    Blue = 8'h26;
end 13'h126f:    begin Red = 8'h60;    Green = 8'h51;    Blue = 8'h30;
end 13'h1270:    begin Red = 8'h69;    Green = 8'h51;    Blue = 8'h39;
end 13'h1271:    begin Red = 8'h57;    Green = 8'h47;    Blue = 8'h38;
end 13'h1272:    begin Red = 8'h54;    Green = 8'h49;    Blue = 8'h2b;
end 13'h1273:    begin Red = 8'hf4;    Green = 8'hd1;    Blue = 8'hab;
end 13'h1274:    begin Red = 8'ha4;    Green = 8'h99;    Blue = 8'h7b;
end 13'h1275:    begin Red = 8'h81;    Green = 8'h66;    Blue = 8'h55;
end 13'h1276:    begin Red = 8'h73;    Green = 8'h5f;    Blue = 8'h44;
end 13'h1277:    begin Red = 8'h70;    Green = 8'h50;    Blue = 8'h1f;
end 13'h1278:    begin Red = 8'h5e;    Green = 8'h47;    Blue = 8'h25;
end 13'h1279:    begin Red = 8'hfe;    Green = 8'hf2;    Blue = 8'hbe;
end 13'h127a:    begin Red = 8'h87;    Green = 8'h6d;    Blue = 8'h54;
end 13'h127b:    begin Red = 8'h51;    Green = 8'h43;    Blue = 8'h36;
end 13'h127c:    begin Red = 8'h50;    Green = 8'h43;    Blue = 8'h3a;
end 13'h127d:    begin Red = 8'h66;    Green = 8'h4d;    Blue = 8'h46;
end 13'h127e:    begin Red = 8'h62;    Green = 8'h4b;    Blue = 8'h2b;
end 13'h127f:    begin Red = 8'h64;    Green = 8'h4e;    Blue = 8'h29;
end 13'h1280:    begin Red = 8'h5f;    Green = 8'h4b;    Blue = 8'h32;
end 13'h1281:    begin Red = 8'h6a;    Green = 8'h57;    Blue = 8'h50;
end 13'h1282:    begin Red = 8'hc4;    Green = 8'hc4;    Blue = 8'hb1;
end 13'h1283:    begin Red = 8'hc7;    Green = 8'ha4;    Blue = 8'h5a;
end 13'h1284:    begin Red = 8'hc1;    Green = 8'ha5;    Blue = 8'h65;
end 13'h1285:    begin Red = 8'hce;    Green = 8'ha7;    Blue = 8'h69;
end 13'h1286:    begin Red = 8'hd2;    Green = 8'hb2;    Blue = 8'h72;
end 13'h1287:    begin Red = 8'hd9;    Green = 8'hd0;    Blue = 8'hc0;
end 13'h1288:    begin Red = 8'hbe;    Green = 8'ha5;    Blue = 8'h7d;
end 13'h1289:    begin Red = 8'hd1;    Green = 8'hb6;    Blue = 8'h98;
end 13'h128a:    begin Red = 8'h46;    Green = 8'h3b;    Blue = 8'h39;
end 13'h128b:    begin Red = 8'h36;    Green = 8'h34;    Blue = 8'h34;
end 13'h128c:    begin Red = 8'he5;    Green = 8'hc2;    Blue = 8'h9c;
end 13'h128d:    begin Red = 8'hee;    Green = 8'hc8;    Blue = 8'ha1;
end 13'h128e:    begin Red = 8'h50;    Green = 8'h3e;    Blue = 8'h28;
end 13'h128f:    begin Red = 8'h5f;    Green = 8'h55;    Blue = 8'h31;
end 13'h1290:    begin Red = 8'h65;    Green = 8'h4b;    Blue = 8'h30;
end 13'h1291:    begin Red = 8'ha4;    Green = 8'h92;    Blue = 8'h6c;
end 13'h1292:    begin Red = 8'h65;    Green = 8'h52;    Blue = 8'h41;
end 13'h1293:    begin Red = 8'h7f;    Green = 8'h64;    Blue = 8'h53;
end 13'h1294:    begin Red = 8'h6c;    Green = 8'h50;    Blue = 8'h2b;
end 13'h1295:    begin Red = 8'h60;    Green = 8'h46;    Blue = 8'h2d;
end 13'h1296:    begin Red = 8'h62;    Green = 8'h4c;    Blue = 8'h27;
end 13'h1297:    begin Red = 8'hfb;    Green = 8'hef;    Blue = 8'hbf;
end 13'h1298:    begin Red = 8'h5e;    Green = 8'h50;    Blue = 8'h36;
end 13'h1299:    begin Red = 8'h60;    Green = 8'h51;    Blue = 8'h3c;
end 13'h129a:    begin Red = 8'h4c;    Green = 8'h45;    Blue = 8'h2b;
end 13'h129b:    begin Red = 8'h61;    Green = 8'h4f;    Blue = 8'h45;
end 13'h129c:    begin Red = 8'h65;    Green = 8'h4d;    Blue = 8'h35;
end 13'h129d:    begin Red = 8'h97;    Green = 8'h91;    Blue = 8'h84;
end 13'h129e:    begin Red = 8'hc0;    Green = 8'ha0;    Blue = 8'h58;
end 13'h129f:    begin Red = 8'hc7;    Green = 8'hab;    Blue = 8'h6c;
end 13'h12a0:    begin Red = 8'hb6;    Green = 8'h9b;    Blue = 8'h61;
end 13'h12a1:    begin Red = 8'hc4;    Green = 8'h9f;    Blue = 8'h5f;
end 13'h12a2:    begin Red = 8'h46;    Green = 8'h3f;    Blue = 8'h35;
end 13'h12a3:    begin Red = 8'h40;    Green = 8'h40;    Blue = 8'h36;
end 13'h12a4:    begin Red = 8'hc5;    Green = 8'hae;    Blue = 8'h93;
end 13'h12a5:    begin Red = 8'hb0;    Green = 8'h94;    Blue = 8'h73;
end 13'h12a6:    begin Red = 8'hcc;    Green = 8'hc3;    Blue = 8'h9f;
end 13'h12a7:    begin Red = 8'h53;    Green = 8'h4a;    Blue = 8'h3b;
end 13'h12a8:    begin Red = 8'h4c;    Green = 8'h3b;    Blue = 8'h27;
end 13'h12a9:    begin Red = 8'h63;    Green = 8'h4a;    Blue = 8'h34;
end 13'h12aa:    begin Red = 8'h4e;    Green = 8'h3a;    Blue = 8'h21;
end 13'h12ab:    begin Red = 8'hed;    Green = 8'hd5;    Blue = 8'ha5;
end 13'h12ac:    begin Red = 8'h56;    Green = 8'h54;    Blue = 8'h45;
end 13'h12ad:    begin Red = 8'h7c;    Green = 8'h61;    Blue = 8'h34;
end 13'h12ae:    begin Red = 8'h57;    Green = 8'h52;    Blue = 8'h4c;
end 13'h12af:    begin Red = 8'h73;    Green = 8'h54;    Blue = 8'h28;
end 13'h12b0:    begin Red = 8'h62;    Green = 8'h4d;    Blue = 8'h52;
end 13'h12b1:    begin Red = 8'h03;    Green = 8'hb2;    Blue = 8'h80;
end 13'h12b2:    begin Red = 8'h46;    Green = 8'h3f;    Blue = 8'h23;
end 13'h12b3:    begin Red = 8'h5b;    Green = 8'h46;    Blue = 8'h35;
end 13'h12b4:    begin Red = 8'h56;    Green = 8'h46;    Blue = 8'h2d;
end 13'h12b5:    begin Red = 8'h4a;    Green = 8'h38;    Blue = 8'h2a;
end 13'h12b6:    begin Red = 8'h2e;    Green = 8'h1d;    Blue = 8'h13;
end 13'h12b7:    begin Red = 8'h56;    Green = 8'h3c;    Blue = 8'h2b;
end 13'h12b8:    begin Red = 8'h5a;    Green = 8'h39;    Blue = 8'h26;
end 13'h12b9:    begin Red = 8'h52;    Green = 8'h37;    Blue = 8'h2c;
end 13'h12ba:    begin Red = 8'h4e;    Green = 8'h42;    Blue = 8'h2c;
end 13'h12bb:    begin Red = 8'ha9;    Green = 8'h90;    Blue = 8'h80;
end 13'h12bc:    begin Red = 8'ha5;    Green = 8'h8c;    Blue = 8'h4b;
end 13'h12bd:    begin Red = 8'hb7;    Green = 8'ha0;    Blue = 8'h68;
end 13'h12be:    begin Red = 8'hc3;    Green = 8'ha2;    Blue = 8'h62;
end 13'h12bf:    begin Red = 8'hb1;    Green = 8'h99;    Blue = 8'h5f;
end 13'h12c0:    begin Red = 8'hb6;    Green = 8'h9c;    Blue = 8'h6d;
end 13'h12c1:    begin Red = 8'hd2;    Green = 8'hd0;    Blue = 8'hc4;
end 13'h12c2:    begin Red = 8'hcc;    Green = 8'hc3;    Blue = 8'hac;
end 13'h12c3:    begin Red = 8'h8a;    Green = 8'h83;    Blue = 8'h6a;
end 13'h12c4:    begin Red = 8'hc3;    Green = 8'h8f;    Blue = 8'h55;
end 13'h12c5:    begin Red = 8'hc3;    Green = 8'h92;    Blue = 8'h57;
end 13'h12c6:    begin Red = 8'hc2;    Green = 8'h94;    Blue = 8'h59;
end 13'h12c7:    begin Red = 8'hc5;    Green = 8'h98;    Blue = 8'h5d;
end 13'h12c8:    begin Red = 8'hbd;    Green = 8'h99;    Blue = 8'h5d;
end 13'h12c9:    begin Red = 8'had;    Green = 8'h7e;    Blue = 8'h4a;
end 13'h12ca:    begin Red = 8'hb3;    Green = 8'h88;    Blue = 8'h44;
end 13'h12cb:    begin Red = 8'hb7;    Green = 8'h90;    Blue = 8'h55;
end 13'h12cc:    begin Red = 8'hbe;    Green = 8'h8c;    Blue = 8'h59;
end 13'h12cd:    begin Red = 8'haf;    Green = 8'h89;    Blue = 8'h4b;
end 13'h12ce:    begin Red = 8'hb2;    Green = 8'h89;    Blue = 8'h49;
end 13'h12cf:    begin Red = 8'hb7;    Green = 8'h8e;    Blue = 8'h50;
end 13'h12d0:    begin Red = 8'ha9;    Green = 8'h81;    Blue = 8'h4e;
end 13'h12d1:    begin Red = 8'h90;    Green = 8'h6a;    Blue = 8'h3b;
end 13'h12d2:    begin Red = 8'h95;    Green = 8'h6e;    Blue = 8'h43;
end 13'h12d3:    begin Red = 8'h8e;    Green = 8'h6c;    Blue = 8'h3c;
end 13'h12d4:    begin Red = 8'h81;    Green = 8'h5f;    Blue = 8'h39;
end 13'h12d5:    begin Red = 8'he5;    Green = 8'hd6;    Blue = 8'hcd;
end 13'h12d6:    begin Red = 8'hc8;    Green = 8'hc2;    Blue = 8'h9d;
end 13'h12d7:    begin Red = 8'ha7;    Green = 8'ha3;    Blue = 8'h86;
end 13'h12d8:    begin Red = 8'h46;    Green = 8'h38;    Blue = 8'h1b;
end 13'h12d9:    begin Red = 8'h43;    Green = 8'h33;    Blue = 8'h1a;
end 13'h12da:    begin Red = 8'h5f;    Green = 8'h4c;    Blue = 8'h2c;
end 13'h12db:    begin Red = 8'h4a;    Green = 8'h35;    Blue = 8'h1a;
end 13'h12dc:    begin Red = 8'h50;    Green = 8'h41;    Blue = 8'h2a;
end 13'h12dd:    begin Red = 8'h5d;    Green = 8'h4f;    Blue = 8'h42;
end 13'h12de:    begin Red = 8'h4f;    Green = 8'h3f;    Blue = 8'h25;
end 13'h12df:    begin Red = 8'h80;    Green = 8'h66;    Blue = 8'h4b;
end 13'h12e0:    begin Red = 8'h5d;    Green = 8'h4a;    Blue = 8'h50;
end 13'h12e1:    begin Red = 8'h7f;    Green = 8'h5e;    Blue = 8'h28;
end 13'h12e2:    begin Red = 8'h6d;    Green = 8'h56;    Blue = 8'h22;
end 13'h12e3:    begin Red = 8'h59;    Green = 8'h47;    Blue = 8'h17;
end 13'h12e4:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h95;
end 13'h12e5:    begin Red = 8'h5c;    Green = 8'h50;    Blue = 8'h3a;
end 13'h12e6:    begin Red = 8'h59;    Green = 8'h4a;    Blue = 8'h35;
end 13'h12e7:    begin Red = 8'h54;    Green = 8'h46;    Blue = 8'h23;
end 13'h12e8:    begin Red = 8'h48;    Green = 8'h34;    Blue = 8'h2b;
end 13'h12e9:    begin Red = 8'h68;    Green = 8'h59;    Blue = 8'h44;
end 13'h12ea:    begin Red = 8'h02;    Green = 8'hf1;    Blue = 8'hff;
end 13'h12eb:    begin Red = 8'h4a;    Green = 8'h3e;    Blue = 8'h26;
end 13'h12ec:    begin Red = 8'h04;    Green = 8'hf2;    Blue = 8'hf6;
end 13'h12ed:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'hdb;
end 13'h12ee:    begin Red = 8'h43;    Green = 8'h30;    Blue = 8'h10;
end 13'h12ef:    begin Red = 8'h49;    Green = 8'h42;    Blue = 8'h28;
end 13'h12f0:    begin Red = 8'h53;    Green = 8'h3a;    Blue = 8'h33;
end 13'h12f1:    begin Red = 8'hab;    Green = 8'h8e;    Blue = 8'h7b;
end 13'h12f2:    begin Red = 8'h9b;    Green = 8'h7a;    Blue = 8'h6f;
end 13'h12f3:    begin Red = 8'h9b;    Green = 8'h7e;    Blue = 8'h70;
end 13'h12f4:    begin Red = 8'h9f;    Green = 8'h87;    Blue = 8'h4f;
end 13'h12f5:    begin Red = 8'hbe;    Green = 8'ha0;    Blue = 8'h65;
end 13'h12f6:    begin Red = 8'hc0;    Green = 8'ha0;    Blue = 8'h60;
end 13'h12f7:    begin Red = 8'hb2;    Green = 8'h96;    Blue = 8'h60;
end 13'h12f8:    begin Red = 8'hc7;    Green = 8'hc7;    Blue = 8'hb8;
end 13'h12f9:    begin Red = 8'he2;    Green = 8'hdd;    Blue = 8'hc3;
end 13'h12fa:    begin Red = 8'h8f;    Green = 8'h8a;    Blue = 8'h75;
end 13'h12fb:    begin Red = 8'h76;    Green = 8'h5d;    Blue = 8'h39;
end 13'h12fc:    begin Red = 8'h6c;    Green = 8'h58;    Blue = 8'h38;
end 13'h12fd:    begin Red = 8'h6f;    Green = 8'h58;    Blue = 8'h3d;
end 13'h12fe:    begin Red = 8'h72;    Green = 8'h65;    Blue = 8'h5b;
end 13'h12ff:    begin Red = 8'hdd;    Green = 8'hd7;    Blue = 8'hc0;
end 13'h1300:    begin Red = 8'hbe;    Green = 8'h8b;    Blue = 8'h54;
end 13'h1301:    begin Red = 8'hb8;    Green = 8'h8b;    Blue = 8'h52;
end 13'h1302:    begin Red = 8'hb2;    Green = 8'h8c;    Blue = 8'h4e;
end 13'h1303:    begin Red = 8'hbc;    Green = 8'h8b;    Blue = 8'h50;
end 13'h1304:    begin Red = 8'hbc;    Green = 8'h88;    Blue = 8'h4e;
end 13'h1305:    begin Red = 8'hb5;    Green = 8'h87;    Blue = 8'h4c;
end 13'h1306:    begin Red = 8'hbe;    Green = 8'h93;    Blue = 8'h44;
end 13'h1307:    begin Red = 8'hb4;    Green = 8'h8c;    Blue = 8'h51;
end 13'h1308:    begin Red = 8'hb1;    Green = 8'h86;    Blue = 8'h51;
end 13'h1309:    begin Red = 8'hac;    Green = 8'h84;    Blue = 8'h47;
end 13'h130a:    begin Red = 8'ha9;    Green = 8'h81;    Blue = 8'h43;
end 13'h130b:    begin Red = 8'h84;    Green = 8'h60;    Blue = 8'h30;
end 13'h130c:    begin Red = 8'h8d;    Green = 8'h68;    Blue = 8'h3b;
end 13'h130d:    begin Red = 8'h88;    Green = 8'h69;    Blue = 8'h32;
end 13'h130e:    begin Red = 8'h86;    Green = 8'h6a;    Blue = 8'h3a;
end 13'h130f:    begin Red = 8'h8a;    Green = 8'h64;    Blue = 8'h33;
end 13'h1310:    begin Red = 8'h77;    Green = 8'h5a;    Blue = 8'h2e;
end 13'h1311:    begin Red = 8'h55;    Green = 8'h4a;    Blue = 8'h38;
end 13'h1312:    begin Red = 8'h2f;    Green = 8'h27;    Blue = 8'h1a;
end 13'h1313:    begin Red = 8'hfc;    Green = 8'hf6;    Blue = 8'hc2;
end 13'h1314:    begin Red = 8'h02;    Green = 8'hc1;    Blue = 8'hbb;
end 13'h1315:    begin Red = 8'h54;    Green = 8'h3e;    Blue = 8'h27;
end 13'h1316:    begin Red = 8'h6a;    Green = 8'h82;    Blue = 8'ha4;
end 13'h1317:    begin Red = 8'h6f;    Green = 8'h84;    Blue = 8'hbb;
end 13'h1318:    begin Red = 8'h56;    Green = 8'h3d;    Blue = 8'h1f;
end 13'h1319:    begin Red = 8'hab;    Green = 8'ha8;    Blue = 8'h9c;
end 13'h131a:    begin Red = 8'haa;    Green = 8'h8c;    Blue = 8'h58;
end 13'h131b:    begin Red = 8'hd8;    Green = 8'hcf;    Blue = 8'hb9;
end 13'h131c:    begin Red = 8'hff;    Green = 8'hfe;    Blue = 8'he2;
end 13'h131d:    begin Red = 8'h55;    Green = 8'h4e;    Blue = 8'h4f;
end 13'h131e:    begin Red = 8'h8c;    Green = 8'hab;    Blue = 8'hd9;
end 13'h131f:    begin Red = 8'h8c;    Green = 8'h9c;    Blue = 8'hbe;
end 13'h1320:    begin Red = 8'h93;    Green = 8'ha9;    Blue = 8'hdb;
end 13'h1321:    begin Red = 8'hd7;    Green = 8'hab;    Blue = 8'h6e;
end 13'h1322:    begin Red = 8'hee;    Green = 8'hc5;    Blue = 8'h83;
end 13'h1323:    begin Red = 8'he9;    Green = 8'hc2;    Blue = 8'h7f;
end 13'h1324:    begin Red = 8'he9;    Green = 8'hbf;    Blue = 8'h83;
end 13'h1325:    begin Red = 8'hda;    Green = 8'hac;    Blue = 8'h70;
end 13'h1326:    begin Red = 8'hc3;    Green = 8'h9c;    Blue = 8'h63;
end 13'h1327:    begin Red = 8'he5;    Green = 8'he8;    Blue = 8'hd7;
end 13'h1328:    begin Red = 8'hd0;    Green = 8'ha4;    Blue = 8'h63;
end 13'h1329:    begin Red = 8'hd3;    Green = 8'ha7;    Blue = 8'h6a;
end 13'h132a:    begin Red = 8'he2;    Green = 8'hbb;    Blue = 8'h7a;
end 13'h132b:    begin Red = 8'hdf;    Green = 8'hba;    Blue = 8'h76;
end 13'h132c:    begin Red = 8'hde;    Green = 8'hb5;    Blue = 8'h75;
end 13'h132d:    begin Red = 8'hcb;    Green = 8'h9f;    Blue = 8'h62;
end 13'h132e:    begin Red = 8'hb9;    Green = 8'h8d;    Blue = 8'h5e;
end 13'h132f:    begin Red = 8'ha0;    Green = 8'h82;    Blue = 8'h5b;
end 13'h1330:    begin Red = 8'hab;    Green = 8'h8f;    Blue = 8'h6d;
end 13'h1331:    begin Red = 8'hcc;    Green = 8'ha6;    Blue = 8'h7f;
end 13'h1332:    begin Red = 8'hb7;    Green = 8'h92;    Blue = 8'h5e;
end 13'h1333:    begin Red = 8'hb5;    Green = 8'h8f;    Blue = 8'h5e;
end 13'h1334:    begin Red = 8'hb0;    Green = 8'h91;    Blue = 8'h5a;
end 13'h1335:    begin Red = 8'hb3;    Green = 8'h97;    Blue = 8'h58;
end 13'h1336:    begin Red = 8'ha0;    Green = 8'h7a;    Blue = 8'h4b;
end 13'h1337:    begin Red = 8'h8c;    Green = 8'h6a;    Blue = 8'h3d;
end 13'h1338:    begin Red = 8'h8f;    Green = 8'h6f;    Blue = 8'h46;
end 13'h1339:    begin Red = 8'hee;    Green = 8'hd5;    Blue = 8'had;
end 13'h133a:    begin Red = 8'he8;    Green = 8'hc6;    Blue = 8'ha3;
end 13'h133b:    begin Red = 8'hf0;    Green = 8'hd6;    Blue = 8'ha3;
end 13'h133c:    begin Red = 8'h96;    Green = 8'h80;    Blue = 8'h5b;
end 13'h133d:    begin Red = 8'h99;    Green = 8'h87;    Blue = 8'h63;
end 13'h133e:    begin Red = 8'hec;    Green = 8'hc8;    Blue = 8'h98;
end 13'h133f:    begin Red = 8'hf9;    Green = 8'hd7;    Blue = 8'haa;
end 13'h1340:    begin Red = 8'he2;    Green = 8'hc3;    Blue = 8'h95;
end 13'h1341:    begin Red = 8'h46;    Green = 8'h46;    Blue = 8'h20;
end 13'h1342:    begin Red = 8'h50;    Green = 8'h3d;    Blue = 8'h1f;
end 13'h1343:    begin Red = 8'hba;    Green = 8'h9c;    Blue = 8'h65;
end 13'h1344:    begin Red = 8'hca;    Green = 8'hae;    Blue = 8'h71;
end 13'h1345:    begin Red = 8'hce;    Green = 8'hac;    Blue = 8'h70;
end 13'h1346:    begin Red = 8'hde;    Green = 8'hd5;    Blue = 8'hc2;
end 13'h1347:    begin Red = 8'h5d;    Green = 8'h51;    Blue = 8'h4d;
end 13'h1348:    begin Red = 8'hd4;    Green = 8'had;    Blue = 8'h6c;
end 13'h1349:    begin Red = 8'h06;    Green = 8'h93;    Blue = 8'hc0;
end 13'h134a:    begin Red = 8'h08;    Green = 8'h14;    Blue = 8'hf8;
end 13'h134b:    begin Red = 8'h07;    Green = 8'hf5;    Blue = 8'h08;
end 13'h134c:    begin Red = 8'h07;    Green = 8'hf4;    Blue = 8'heb;
end 13'h134d:    begin Red = 8'h06;    Green = 8'h94;    Blue = 8'h13;
end 13'h134e:    begin Red = 8'h05;    Green = 8'h02;    Blue = 8'hb0;
end 13'h134f:    begin Red = 8'h8a;    Green = 8'h63;    Blue = 8'h3a;
end 13'h1350:    begin Red = 8'h8d;    Green = 8'h73;    Blue = 8'h42;
end 13'h1351:    begin Red = 8'hcf;    Green = 8'ha6;    Blue = 8'h6e;
end 13'h1352:    begin Red = 8'hc7;    Green = 8'h9e;    Blue = 8'h66;
end 13'h1353:    begin Red = 8'hc9;    Green = 8'ha1;    Blue = 8'h6d;
end 13'h1354:    begin Red = 8'hca;    Green = 8'h9f;    Blue = 8'h68;
end 13'h1355:    begin Red = 8'hc6;    Green = 8'h9e;    Blue = 8'h6a;
end 13'h1356:    begin Red = 8'hc8;    Green = 8'h9b;    Blue = 8'h64;
end 13'h1357:    begin Red = 8'hc2;    Green = 8'h9b;    Blue = 8'h60;
end 13'h1358:    begin Red = 8'hd0;    Green = 8'ha8;    Blue = 8'h62;
end 13'h1359:    begin Red = 8'hd2;    Green = 8'ha4;    Blue = 8'h66;
end 13'h135a:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'ha0;
end 13'h135b:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'heb;
end 13'h135c:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'hc8;
end 13'h135d:    begin Red = 8'h07;    Green = 8'h94;    Blue = 8'hc9;
end 13'h135e:    begin Red = 8'h07;    Green = 8'h44;    Blue = 8'hed;
end 13'h135f:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'hc5;
end 13'h1360:    begin Red = 8'h05;    Green = 8'h22;    Blue = 8'h42;
end 13'h1361:    begin Red = 8'hb3;    Green = 8'h8f;    Blue = 8'h55;
end 13'h1362:    begin Red = 8'h8e;    Green = 8'h63;    Blue = 8'h40;
end 13'h1363:    begin Red = 8'hbd;    Green = 8'h96;    Blue = 8'h5f;
end 13'h1364:    begin Red = 8'hb5;    Green = 8'h8e;    Blue = 8'h57;
end 13'h1365:    begin Red = 8'hdd;    Green = 8'he5;    Blue = 8'hca;
end 13'h1366:    begin Red = 8'ha4;    Green = 8'h83;    Blue = 8'h4e;
end 13'h1367:    begin Red = 8'h06;    Green = 8'h23;    Blue = 8'hea;
end 13'h1368:    begin Red = 8'h06;    Green = 8'h23;    Blue = 8'hf7;
end 13'h1369:    begin Red = 8'h06;    Green = 8'h13;    Blue = 8'hc5;
end 13'h136a:    begin Red = 8'h05;    Green = 8'he3;    Blue = 8'hd8;
end 13'h136b:    begin Red = 8'h05;    Green = 8'hd3;    Blue = 8'hf3;
end 13'h136c:    begin Red = 8'h04;    Green = 8'hb3;    Blue = 8'h05;
end 13'h136d:    begin Red = 8'hf4;    Green = 8'hdc;    Blue = 8'hae;
end 13'h136e:    begin Red = 8'haa;    Green = 8'h97;    Blue = 8'h6f;
end 13'h136f:    begin Red = 8'hb3;    Green = 8'h95;    Blue = 8'h71;
end 13'h1370:    begin Red = 8'hea;    Green = 8'hc4;    Blue = 8'h97;
end 13'h1371:    begin Red = 8'heb;    Green = 8'hcb;    Blue = 8'h9c;
end 13'h1372:    begin Red = 8'he5;    Green = 8'hc3;    Blue = 8'h93;
end 13'h1373:    begin Red = 8'h9e;    Green = 8'h81;    Blue = 8'h61;
end 13'h1374:    begin Red = 8'he3;    Green = 8'hc9;    Blue = 8'h98;
end 13'h1375:    begin Red = 8'he1;    Green = 8'hc7;    Blue = 8'h94;
end 13'h1376:    begin Red = 8'h02;    Green = 8'he1;    Blue = 8'h8b;
end 13'h1377:    begin Red = 8'h59;    Green = 8'h3e;    Blue = 8'h2d;
end 13'h1378:    begin Red = 8'hbd;    Green = 8'h9c;    Blue = 8'h53;
end 13'h1379:    begin Red = 8'hc3;    Green = 8'ha1;    Blue = 8'h5d;
end 13'h137a:    begin Red = 8'he2;    Green = 8'hdb;    Blue = 8'hc9;
end 13'h137b:    begin Red = 8'h52;    Green = 8'h4d;    Blue = 8'h48;
end 13'h137c:    begin Red = 8'h42;    Green = 8'h3e;    Blue = 8'h3f;
end 13'h137d:    begin Red = 8'hd6;    Green = 8'ha9;    Blue = 8'h68;
end 13'h137e:    begin Red = 8'h06;    Green = 8'hc3;    Blue = 8'hc0;
end 13'h137f:    begin Red = 8'h07;    Green = 8'hc4;    Blue = 8'hfb;
end 13'h1380:    begin Red = 8'h08;    Green = 8'h05;    Blue = 8'h1d;
end 13'h1381:    begin Red = 8'h08;    Green = 8'h45;    Blue = 8'h05;
end 13'h1382:    begin Red = 8'h08;    Green = 8'h24;    Blue = 8'hfe;
end 13'h1383:    begin Red = 8'h06;    Green = 8'h64;    Blue = 8'h1a;
end 13'h1384:    begin Red = 8'h05;    Green = 8'h72;    Blue = 8'hb6;
end 13'h1385:    begin Red = 8'h91;    Green = 8'h6f;    Blue = 8'h3f;
end 13'h1386:    begin Red = 8'ha9;    Green = 8'h84;    Blue = 8'h50;
end 13'h1387:    begin Red = 8'hc5;    Green = 8'h9a;    Blue = 8'h67;
end 13'h1388:    begin Red = 8'hd4;    Green = 8'ha9;    Blue = 8'h65;
end 13'h1389:    begin Red = 8'hce;    Green = 8'ha1;    Blue = 8'h68;
end 13'h138a:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'h80;
end 13'h138b:    begin Red = 8'h07;    Green = 8'hb5;    Blue = 8'h17;
end 13'h138c:    begin Red = 8'h07;    Green = 8'hd4;    Blue = 8'hbc;
end 13'h138d:    begin Red = 8'h07;    Green = 8'h64;    Blue = 8'he9;
end 13'h138e:    begin Red = 8'h07;    Green = 8'h85;    Blue = 8'h08;
end 13'h138f:    begin Red = 8'h06;    Green = 8'h43;    Blue = 8'h9c;
end 13'h1390:    begin Red = 8'h05;    Green = 8'h32;    Blue = 8'he4;
end 13'h1391:    begin Red = 8'hb8;    Green = 8'h95;    Blue = 8'h5d;
end 13'h1392:    begin Red = 8'hb6;    Green = 8'h8e;    Blue = 8'h5b;
end 13'h1393:    begin Red = 8'ha3;    Green = 8'h7e;    Blue = 8'h51;
end 13'h1394:    begin Red = 8'h06;    Green = 8'h44;    Blue = 8'h3d;
end 13'h1395:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'hd7;
end 13'h1396:    begin Red = 8'h06;    Green = 8'h13;    Blue = 8'hd9;
end 13'h1397:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'hca;
end 13'h1398:    begin Red = 8'h04;    Green = 8'hd2;    Blue = 8'he2;
end 13'h1399:    begin Red = 8'h8d;    Green = 8'h6a;    Blue = 8'h44;
end 13'h139a:    begin Red = 8'hdf;    Green = 8'hd6;    Blue = 8'hae;
end 13'h139b:    begin Red = 8'hc0;    Green = 8'hc7;    Blue = 8'ha5;
end 13'h139c:    begin Red = 8'h65;    Green = 8'h4c;    Blue = 8'h4f;
end 13'h139d:    begin Red = 8'h62;    Green = 8'h4d;    Blue = 8'h4a;
end 13'h139e:    begin Red = 8'h8f;    Green = 8'h70;    Blue = 8'h6d;
end 13'h139f:    begin Red = 8'h8d;    Green = 8'h6b;    Blue = 8'h6a;
end 13'h13a0:    begin Red = 8'h8b;    Green = 8'h69;    Blue = 8'h68;
end 13'h13a1:    begin Red = 8'h70;    Green = 8'h54;    Blue = 8'h53;
end 13'h13a2:    begin Red = 8'h73;    Green = 8'h59;    Blue = 8'h58;
end 13'h13a3:    begin Red = 8'h8c;    Green = 8'h6c;    Blue = 8'h6d;
end 13'h13a4:    begin Red = 8'h75;    Green = 8'h5b;    Blue = 8'h5a;
end 13'h13a5:    begin Red = 8'h8e;    Green = 8'h6b;    Blue = 8'h71;
end 13'h13a6:    begin Red = 8'h8a;    Green = 8'h69;    Blue = 8'h64;
end 13'h13a7:    begin Red = 8'h58;    Green = 8'h3e;    Blue = 8'h4b;
end 13'h13a8:    begin Red = 8'h7a;    Green = 8'h57;    Blue = 8'h5d;
end 13'h13a9:    begin Red = 8'h97;    Green = 8'h6f;    Blue = 8'h70;
end 13'h13aa:    begin Red = 8'h8a;    Green = 8'h6a;    Blue = 8'h6b;
end 13'h13ab:    begin Red = 8'h75;    Green = 8'h56;    Blue = 8'h5b;
end 13'h13ac:    begin Red = 8'h5c;    Green = 8'h3a;    Blue = 8'h48;
end 13'h13ad:    begin Red = 8'h8e;    Green = 8'h61;    Blue = 8'h64;
end 13'h13ae:    begin Red = 8'h79;    Green = 8'h5d;    Blue = 8'h5c;
end 13'h13af:    begin Red = 8'h92;    Green = 8'h70;    Blue = 8'h71;
end 13'h13b0:    begin Red = 8'h6c;    Green = 8'h54;    Blue = 8'h52;
end 13'h13b1:    begin Red = 8'h5f;    Green = 8'h41;    Blue = 8'h4d;
end 13'h13b2:    begin Red = 8'hf3;    Green = 8'hd4;    Blue = 8'ha5;
end 13'h13b3:    begin Red = 8'hff;    Green = 8'hf1;    Blue = 8'hd0;
end 13'h13b4:    begin Red = 8'hfa;    Green = 8'hdd;    Blue = 8'hb5;
end 13'h13b5:    begin Red = 8'h4d;    Green = 8'h48;    Blue = 8'h3f;
end 13'h13b6:    begin Red = 8'h55;    Green = 8'h52;    Blue = 8'h49;
end 13'h13b7:    begin Red = 8'hc3;    Green = 8'hb9;    Blue = 8'ha7;
end 13'h13b8:    begin Red = 8'h90;    Green = 8'h93;    Blue = 8'h7a;
end 13'h13b9:    begin Red = 8'hee;    Green = 8'hc4;    Blue = 8'h8a;
end 13'h13ba:    begin Red = 8'h8b;    Green = 8'h56;    Blue = 8'h14;
end 13'h13bb:    begin Red = 8'h06;    Green = 8'hc4;    Blue = 8'h54;
end 13'h13bc:    begin Red = 8'hd7;    Green = 8'hae;    Blue = 8'h70;
end 13'h13bd:    begin Red = 8'h7b;    Green = 8'h5b;    Blue = 8'h32;
end 13'h13be:    begin Red = 8'h85;    Green = 8'h64;    Blue = 8'h37;
end 13'h13bf:    begin Red = 8'hc1;    Green = 8'h98;    Blue = 8'h56;
end 13'h13c0:    begin Red = 8'hbb;    Green = 8'h8e;    Blue = 8'h55;
end 13'h13c1:    begin Red = 8'hbd;    Green = 8'h90;    Blue = 8'h57;
end 13'h13c2:    begin Red = 8'hda;    Green = 8'hae;    Blue = 8'h6d;
end 13'h13c3:    begin Red = 8'hf6;    Green = 8'hd4;    Blue = 8'h97;
end 13'h13c4:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'ha8;
end 13'h13c5:    begin Red = 8'h06;    Green = 8'h23;    Blue = 8'hcd;
end 13'h13c6:    begin Red = 8'hb9;    Green = 8'h92;    Blue = 8'h5b;
end 13'h13c7:    begin Red = 8'h78;    Green = 8'h5d;    Blue = 8'h32;
end 13'h13c8:    begin Red = 8'h8f;    Green = 8'h62;    Blue = 8'h39;
end 13'h13c9:    begin Red = 8'ha6;    Green = 8'h7e;    Blue = 8'h4b;
end 13'h13ca:    begin Red = 8'h9d;    Green = 8'h7d;    Blue = 8'h4c;
end 13'h13cb:    begin Red = 8'ha3;    Green = 8'h74;    Blue = 8'h46;
end 13'h13cc:    begin Red = 8'h98;    Green = 8'h76;    Blue = 8'h46;
end 13'h13cd:    begin Red = 8'h8f;    Green = 8'h6b;    Blue = 8'h49;
end 13'h13ce:    begin Red = 8'ha7;    Green = 8'h83;    Blue = 8'h53;
end 13'h13cf:    begin Red = 8'h05;    Green = 8'he3;    Blue = 8'ha8;
end 13'h13d0:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'hf5;
end 13'h13d1:    begin Red = 8'h03;    Green = 8'hf2;    Blue = 8'h10;
end 13'h13d2:    begin Red = 8'h78;    Green = 8'h5f;    Blue = 8'h62;
end 13'h13d3:    begin Red = 8'h71;    Green = 8'h57;    Blue = 8'h56;
end 13'h13d4:    begin Red = 8'ha5;    Green = 8'h7d;    Blue = 8'h7e;
end 13'h13d5:    begin Red = 8'ha6;    Green = 8'h7f;    Blue = 8'h80;
end 13'h13d6:    begin Red = 8'ha9;    Green = 8'h86;    Blue = 8'h84;
end 13'h13d7:    begin Red = 8'hac;    Green = 8'h84;    Blue = 8'h85;
end 13'h13d8:    begin Red = 8'ha2;    Green = 8'h7b;    Blue = 8'h7c;
end 13'h13d9:    begin Red = 8'h87;    Green = 8'h68;    Blue = 8'h66;
end 13'h13da:    begin Red = 8'ha8;    Green = 8'h80;    Blue = 8'h76;
end 13'h13db:    begin Red = 8'h6d;    Green = 8'h52;    Blue = 8'h5b;
end 13'h13dc:    begin Red = 8'ha3;    Green = 8'h81;    Blue = 8'h77;
end 13'h13dd:    begin Red = 8'ha1;    Green = 8'h7f;    Blue = 8'h7e;
end 13'h13de:    begin Red = 8'h85;    Green = 8'h69;    Blue = 8'h68;
end 13'h13df:    begin Red = 8'h73;    Green = 8'h51;    Blue = 8'h62;
end 13'h13e0:    begin Red = 8'hfe;    Green = 8'hf1;    Blue = 8'hc7;
end 13'h13e1:    begin Red = 8'h78;    Green = 8'h5a;    Blue = 8'h64;
end 13'h13e2:    begin Red = 8'hb1;    Green = 8'h87;    Blue = 8'h88;
end 13'h13e3:    begin Red = 8'hac;    Green = 8'h7d;    Blue = 8'h83;
end 13'h13e4:    begin Red = 8'h86;    Green = 8'h6e;    Blue = 8'h6c;
end 13'h13e5:    begin Red = 8'hb0;    Green = 8'h7f;    Blue = 8'h83;
end 13'h13e6:    begin Red = 8'had;    Green = 8'h81;    Blue = 8'h82;
end 13'h13e7:    begin Red = 8'h92;    Green = 8'h6b;    Blue = 8'h6e;
end 13'h13e8:    begin Red = 8'hd4;    Green = 8'hba;    Blue = 8'h7f;
end 13'h13e9:    begin Red = 8'hfa;    Green = 8'he4;    Blue = 8'hbb;
end 13'h13ea:    begin Red = 8'hc5;    Green = 8'ha3;    Blue = 8'h51;
end 13'h13eb:    begin Red = 8'hac;    Green = 8'h8c;    Blue = 8'h4f;
end 13'h13ec:    begin Red = 8'hdb;    Green = 8'hd2;    Blue = 8'hbd;
end 13'h13ed:    begin Red = 8'hbd;    Green = 8'hbb;    Blue = 8'ha9;
end 13'h13ee:    begin Red = 8'hd0;    Green = 8'hc7;    Blue = 8'hb6;
end 13'h13ef:    begin Red = 8'hd9;    Green = 8'hd8;    Blue = 8'hbf;
end 13'h13f0:    begin Red = 8'heb;    Green = 8'hc8;    Blue = 8'h88;
end 13'h13f1:    begin Red = 8'h07;    Green = 8'hd4;    Blue = 8'hca;
end 13'h13f2:    begin Red = 8'h88;    Green = 8'h53;    Blue = 8'h11;
end 13'h13f3:    begin Red = 8'h06;    Green = 8'h74;    Blue = 8'h05;
end 13'h13f4:    begin Red = 8'hd2;    Green = 8'ha9;    Blue = 8'h73;
end 13'h13f5:    begin Red = 8'h64;    Green = 8'h4b;    Blue = 8'h23;
end 13'h13f6:    begin Red = 8'h65;    Green = 8'h47;    Blue = 8'h2b;
end 13'h13f7:    begin Red = 8'h9f;    Green = 8'h78;    Blue = 8'h3f;
end 13'h13f8:    begin Red = 8'h9b;    Green = 8'h71;    Blue = 8'h41;
end 13'h13f9:    begin Red = 8'h97;    Green = 8'h72;    Blue = 8'h3e;
end 13'h13fa:    begin Red = 8'h98;    Green = 8'h71;    Blue = 8'h3a;
end 13'h13fb:    begin Red = 8'h96;    Green = 8'h6e;    Blue = 8'h3b;
end 13'h13fc:    begin Red = 8'he4;    Green = 8'hbc;    Blue = 8'h7f;
end 13'h13fd:    begin Red = 8'hf9;    Green = 8'hd2;    Blue = 8'h9b;
end 13'h13fe:    begin Red = 8'h07;    Green = 8'ha4;    Blue = 8'hb7;
end 13'h13ff:    begin Red = 8'h05;    Green = 8'hc3;    Blue = 8'h93;
end 13'h1400:    begin Red = 8'h06;    Green = 8'h54;    Blue = 8'h17;
end 13'h1401:    begin Red = 8'hc8;    Green = 8'h99;    Blue = 8'h6b;
end 13'h1402:    begin Red = 8'h5f;    Green = 8'h45;    Blue = 8'h20;
end 13'h1403:    begin Red = 8'h61;    Green = 8'h43;    Blue = 8'h1f;
end 13'h1404:    begin Red = 8'h58;    Green = 8'h41;    Blue = 8'h1f;
end 13'h1405:    begin Red = 8'h89;    Green = 8'h6b;    Blue = 8'h39;
end 13'h1406:    begin Red = 8'h83;    Green = 8'h63;    Blue = 8'h34;
end 13'h1407:    begin Red = 8'h7f;    Green = 8'h53;    Blue = 8'h22;
end 13'h1408:    begin Red = 8'h7b;    Green = 8'h59;    Blue = 8'h2c;
end 13'h1409:    begin Red = 8'h7d;    Green = 8'h5a;    Blue = 8'h30;
end 13'h140a:    begin Red = 8'h79;    Green = 8'h57;    Blue = 8'h29;
end 13'h140b:    begin Red = 8'h79;    Green = 8'h54;    Blue = 8'h27;
end 13'h140c:    begin Red = 8'h76;    Green = 8'h56;    Blue = 8'h2f;
end 13'h140d:    begin Red = 8'hcc;    Green = 8'ha5;    Blue = 8'h7a;
end 13'h140e:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'hb6;
end 13'h140f:    begin Red = 8'h03;    Green = 8'h82;    Blue = 8'h00;
end 13'h1410:    begin Red = 8'ha8;    Green = 8'h79;    Blue = 8'h45;
end 13'h1411:    begin Red = 8'h8d;    Green = 8'h6e;    Blue = 8'h40;
end 13'h1412:    begin Red = 8'h82;    Green = 8'h64;    Blue = 8'h62;
end 13'h1413:    begin Red = 8'h9f;    Green = 8'h7c;    Blue = 8'h7a;
end 13'h1414:    begin Red = 8'h73;    Green = 8'h4a;    Blue = 8'h5a;
end 13'h1415:    begin Red = 8'h87;    Green = 8'h65;    Blue = 8'h63;
end 13'h1416:    begin Red = 8'ha2;    Green = 8'h7a;    Blue = 8'h78;
end 13'h1417:    begin Red = 8'haa;    Green = 8'h7e;    Blue = 8'h7d;
end 13'h1418:    begin Red = 8'h89;    Green = 8'h66;    Blue = 8'h6a;
end 13'h1419:    begin Red = 8'h73;    Green = 8'h50;    Blue = 8'h57;
end 13'h141a:    begin Red = 8'h77;    Green = 8'h5a;    Blue = 8'h5c;
end 13'h141b:    begin Red = 8'haa;    Green = 8'h76;    Blue = 8'h82;
end 13'h141c:    begin Red = 8'h81;    Green = 8'h64;    Blue = 8'h66;
end 13'h141d:    begin Red = 8'h8a;    Green = 8'h67;    Blue = 8'h6e;
end 13'h141e:    begin Red = 8'h74;    Green = 8'h4e;    Blue = 8'h59;
end 13'h141f:    begin Red = 8'hec;    Green = 8'hdb;    Blue = 8'ha7;
end 13'h1420:    begin Red = 8'hd4;    Green = 8'hb9;    Blue = 8'h84;
end 13'h1421:    begin Red = 8'hd8;    Green = 8'hbd;    Blue = 8'h86;
end 13'h1422:    begin Red = 8'hf5;    Green = 8'hde;    Blue = 8'haa;
end 13'h1423:    begin Red = 8'hc0;    Green = 8'ha2;    Blue = 8'h55;
end 13'h1424:    begin Red = 8'ha4;    Green = 8'h8d;    Blue = 8'h59;
end 13'h1425:    begin Red = 8'hae;    Green = 8'h91;    Blue = 8'h56;
end 13'h1426:    begin Red = 8'hd3;    Green = 8'hb7;    Blue = 8'h72;
end 13'h1427:    begin Red = 8'hd8;    Green = 8'hd8;    Blue = 8'hc5;
end 13'h1428:    begin Red = 8'h48;    Green = 8'h44;    Blue = 8'h41;
end 13'h1429:    begin Red = 8'hc9;    Green = 8'hca;    Blue = 8'hb9;
end 13'h142a:    begin Red = 8'h08;    Green = 8'h14;    Blue = 8'hed;
end 13'h142b:    begin Red = 8'h08;    Green = 8'h45;    Blue = 8'h2d;
end 13'h142c:    begin Red = 8'h06;    Green = 8'h84;    Blue = 8'h05;
end 13'h142d:    begin Red = 8'h57;    Green = 8'h3f;    Blue = 8'h1d;
end 13'h142e:    begin Red = 8'h6d;    Green = 8'h50;    Blue = 8'h32;
end 13'h142f:    begin Red = 8'h6d;    Green = 8'h4e;    Blue = 8'h22;
end 13'h1430:    begin Red = 8'haa;    Green = 8'h7d;    Blue = 8'h46;
end 13'h1431:    begin Red = 8'ha3;    Green = 8'h74;    Blue = 8'h3c;
end 13'h1432:    begin Red = 8'h9e;    Green = 8'h75;    Blue = 8'h3d;
end 13'h1433:    begin Red = 8'h9d;    Green = 8'h75;    Blue = 8'h41;
end 13'h1434:    begin Red = 8'he4;    Green = 8'hc2;    Blue = 8'h82;
end 13'h1435:    begin Red = 8'hfb;    Green = 8'hd3;    Blue = 8'h96;
end 13'h1436:    begin Red = 8'h05;    Green = 8'hc3;    Blue = 8'hb6;
end 13'h1437:    begin Red = 8'hd2;    Green = 8'ha1;    Blue = 8'h69;
end 13'h1438:    begin Red = 8'hbc;    Green = 8'h94;    Blue = 8'h61;
end 13'h1439:    begin Red = 8'h91;    Green = 8'h72;    Blue = 8'h39;
end 13'h143a:    begin Red = 8'h8b;    Green = 8'h68;    Blue = 8'h30;
end 13'h143b:    begin Red = 8'h8b;    Green = 8'h65;    Blue = 8'h38;
end 13'h143c:    begin Red = 8'hc3;    Green = 8'hd1;    Blue = 8'hb3;
end 13'h143d:    begin Red = 8'h80;    Green = 8'h55;    Blue = 8'h20;
end 13'h143e:    begin Red = 8'h81;    Green = 8'h5f;    Blue = 8'h32;
end 13'h143f:    begin Red = 8'hb5;    Green = 8'h8b;    Blue = 8'h59;
end 13'h1440:    begin Red = 8'hc8;    Green = 8'ha4;    Blue = 8'h74;
end 13'h1441:    begin Red = 8'h05;    Green = 8'h13;    Blue = 8'h05;
end 13'h1442:    begin Red = 8'h03;    Green = 8'hf1;    Blue = 8'hc0;
end 13'h1443:    begin Red = 8'ha8;    Green = 8'h75;    Blue = 8'h7c;
end 13'h1444:    begin Red = 8'h22;    Green = 8'h26;    Blue = 8'h66;
end 13'h1445:    begin Red = 8'h49;    Green = 8'h47;    Blue = 8'h79;
end 13'h1446:    begin Red = 8'h3f;    Green = 8'h47;    Blue = 8'h6c;
end 13'h1447:    begin Red = 8'h43;    Green = 8'h3e;    Blue = 8'h80;
end 13'h1448:    begin Red = 8'h6c;    Green = 8'h70;    Blue = 8'h8e;
end 13'h1449:    begin Red = 8'h67;    Green = 8'h6b;    Blue = 8'h89;
end 13'h144a:    begin Red = 8'h6b;    Green = 8'h6d;    Blue = 8'h89;
end 13'h144b:    begin Red = 8'he5;    Green = 8'he4;    Blue = 8'hd6;
end 13'h144c:    begin Red = 8'hef;    Green = 8'hc6;    Blue = 8'h88;
end 13'h144d:    begin Red = 8'he7;    Green = 8'hbd;    Blue = 8'h81;
end 13'h144e:    begin Red = 8'he7;    Green = 8'hc0;    Blue = 8'h7d;
end 13'h144f:    begin Red = 8'hcc;    Green = 8'h9d;    Blue = 8'h67;
end 13'h1450:    begin Red = 8'hcb;    Green = 8'ha3;    Blue = 8'h65;
end 13'h1451:    begin Red = 8'hb8;    Green = 8'h8d;    Blue = 8'h58;
end 13'h1452:    begin Red = 8'h9b;    Green = 8'h7f;    Blue = 8'h4d;
end 13'h1453:    begin Red = 8'hd4;    Green = 8'hac;    Blue = 8'h7b;
end 13'h1454:    begin Red = 8'hcf;    Green = 8'hab;    Blue = 8'h6d;
end 13'h1455:    begin Red = 8'hd5;    Green = 8'hde;    Blue = 8'hc3;
end 13'h1456:    begin Red = 8'hc4;    Green = 8'h9f;    Blue = 8'h68;
end 13'h1457:    begin Red = 8'hc1;    Green = 8'h9c;    Blue = 8'h68;
end 13'h1458:    begin Red = 8'h78;    Green = 8'h5b;    Blue = 8'h60;
end 13'h1459:    begin Red = 8'h84;    Green = 8'h66;    Blue = 8'h66;
end 13'h145a:    begin Red = 8'ha0;    Green = 8'h77;    Blue = 8'h7b;
end 13'h145b:    begin Red = 8'h9d;    Green = 8'h76;    Blue = 8'h77;
end 13'h145c:    begin Red = 8'ha5;    Green = 8'h81;    Blue = 8'h83;
end 13'h145d:    begin Red = 8'hab;    Green = 8'h7a;    Blue = 8'h7d;
end 13'h145e:    begin Red = 8'ha6;    Green = 8'h79;    Blue = 8'h80;
end 13'h145f:    begin Red = 8'h6c;    Green = 8'h49;    Blue = 8'h4d;
end 13'h1460:    begin Red = 8'h6f;    Green = 8'h50;    Blue = 8'h56;
end 13'h1461:    begin Red = 8'hf7;    Green = 8'hd5;    Blue = 8'haf;
end 13'h1462:    begin Red = 8'hff;    Green = 8'hf2;    Blue = 8'hb5;
end 13'h1463:    begin Red = 8'hb2;    Green = 8'h83;    Blue = 8'h8b;
end 13'h1464:    begin Red = 8'hd3;    Green = 8'hd5;    Blue = 8'haf;
end 13'h1465:    begin Red = 8'ha6;    Green = 8'h73;    Blue = 8'h82;
end 13'h1466:    begin Red = 8'h8b;    Green = 8'h64;    Blue = 8'h67;
end 13'h1467:    begin Red = 8'h84;    Green = 8'h67;    Blue = 8'h61;
end 13'h1468:    begin Red = 8'h74;    Green = 8'h4f;    Blue = 8'h60;
end 13'h1469:    begin Red = 8'h25;    Green = 8'h2b;    Blue = 8'h69;
end 13'h146a:    begin Red = 8'h1e;    Green = 8'h29;    Blue = 8'h61;
end 13'h146b:    begin Red = 8'h1b;    Green = 8'h23;    Blue = 8'h74;
end 13'h146c:    begin Red = 8'ha9;    Green = 8'ha0;    Blue = 8'h9b;
end 13'h146d:    begin Red = 8'ha6;    Green = 8'ha4;    Blue = 8'h9b;
end 13'h146e:    begin Red = 8'ha8;    Green = 8'ha4;    Blue = 8'ha2;
end 13'h146f:    begin Red = 8'ha1;    Green = 8'h96;    Blue = 8'h8c;
end 13'h1470:    begin Red = 8'ha8;    Green = 8'h98;    Blue = 8'h74;
end 13'h1471:    begin Red = 8'hda;    Green = 8'hce;    Blue = 8'hbe;
end 13'h1472:    begin Red = 8'hc8;    Green = 8'hac;    Blue = 8'h69;
end 13'h1473:    begin Red = 8'hbe;    Green = 8'ha0;    Blue = 8'h5d;
end 13'h1474:    begin Red = 8'h4d;    Green = 8'h54;    Blue = 8'h81;
end 13'h1475:    begin Red = 8'h57;    Green = 8'h5d;    Blue = 8'h88;
end 13'h1476:    begin Red = 8'h55;    Green = 8'h5b;    Blue = 8'h80;
end 13'h1477:    begin Red = 8'h7b;    Green = 8'h6c;    Blue = 8'h66;
end 13'h1478:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'h30;
end 13'h1479:    begin Red = 8'h06;    Green = 8'h93;    Blue = 8'h72;
end 13'h147a:    begin Red = 8'h04;    Green = 8'hd2;    Blue = 8'h16;
end 13'h147b:    begin Red = 8'hd4;    Green = 8'ha7;    Blue = 8'h70;
end 13'h147c:    begin Red = 8'ha9;    Green = 8'h7e;    Blue = 8'h5b;
end 13'h147d:    begin Red = 8'hef;    Green = 8'hca;    Blue = 8'h84;
end 13'h147e:    begin Red = 8'he5;    Green = 8'hbe;    Blue = 8'h83;
end 13'h147f:    begin Red = 8'he3;    Green = 8'hbb;    Blue = 8'h76;
end 13'h1480:    begin Red = 8'hca;    Green = 8'ha1;    Blue = 8'h5f;
end 13'h1481:    begin Red = 8'hf3;    Green = 8'hcd;    Blue = 8'h9e;
end 13'h1482:    begin Red = 8'h06;    Green = 8'h13;    Blue = 8'h32;
end 13'h1483:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'h30;
end 13'h1484:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'h37;
end 13'h1485:    begin Red = 8'hd7;    Green = 8'hb3;    Blue = 8'h75;
end 13'h1486:    begin Red = 8'hd1;    Green = 8'haa;    Blue = 8'h6f;
end 13'h1487:    begin Red = 8'hd6;    Green = 8'ha0;    Blue = 8'h60;
end 13'h1488:    begin Red = 8'hbe;    Green = 8'h9b;    Blue = 8'h65;
end 13'h1489:    begin Red = 8'hb8;    Green = 8'h9e;    Blue = 8'h63;
end 13'h148a:    begin Red = 8'hc1;    Green = 8'h9d;    Blue = 8'h7b;
end 13'h148b:    begin Red = 8'h03;    Green = 8'hc1;    Blue = 8'hd1;
end 13'h148c:    begin Red = 8'h00;    Green = 8'h31;    Blue = 8'hf0;
end 13'h148d:    begin Red = 8'h9b;    Green = 8'h74;    Blue = 8'h75;
end 13'h148e:    begin Red = 8'h9c;    Green = 8'h77;    Blue = 8'h7f;
end 13'h148f:    begin Red = 8'ha1;    Green = 8'h78;    Blue = 8'h76;
end 13'h1490:    begin Red = 8'h6f;    Green = 8'h45;    Blue = 8'h59;
end 13'h1491:    begin Red = 8'h8c;    Green = 8'h68;    Blue = 8'h6c;
end 13'h1492:    begin Red = 8'h6d;    Green = 8'h51;    Blue = 8'h4d;
end 13'h1493:    begin Red = 8'h82;    Green = 8'h5c;    Blue = 8'h67;
end 13'h1494:    begin Red = 8'hae;    Green = 8'h7f;    Blue = 8'h79;
end 13'h1495:    begin Red = 8'ha3;    Green = 8'h7b;    Blue = 8'h73;
end 13'h1496:    begin Red = 8'h9d;    Green = 8'ha5;    Blue = 8'h88;
end 13'h1497:    begin Red = 8'ha0;    Green = 8'had;    Blue = 8'h8e;
end 13'h1498:    begin Red = 8'ha3;    Green = 8'h74;    Blue = 8'h7a;
end 13'h1499:    begin Red = 8'h71;    Green = 8'h51;    Blue = 8'h5e;
end 13'h149a:    begin Red = 8'hf8;    Green = 8'hd2;    Blue = 8'ha5;
end 13'h149b:    begin Red = 8'he0;    Green = 8'hb7;    Blue = 8'h99;
end 13'h149c:    begin Red = 8'hfd;    Green = 8'hdc;    Blue = 8'haf;
end 13'h149d:    begin Red = 8'ha8;    Green = 8'ha2;    Blue = 8'h99;
end 13'h149e:    begin Red = 8'h98;    Green = 8'h8b;    Blue = 8'h7e;
end 13'h149f:    begin Red = 8'hbb;    Green = 8'h9a;    Blue = 8'h5f;
end 13'h14a0:    begin Red = 8'hb3;    Green = 8'h9d;    Blue = 8'h63;
end 13'h14a1:    begin Red = 8'hbd;    Green = 8'h9d;    Blue = 8'h6c;
end 13'h14a2:    begin Red = 8'hb3;    Green = 8'h9b;    Blue = 8'h69;
end 13'h14a3:    begin Red = 8'hc7;    Green = 8'hb9;    Blue = 8'hb6;
end 13'h14a4:    begin Red = 8'hcf;    Green = 8'hc3;    Blue = 8'hb3;
end 13'h14a5:    begin Red = 8'hcb;    Green = 8'hbd;    Blue = 8'hac;
end 13'h14a6:    begin Red = 8'he8;    Green = 8'hbf;    Blue = 8'h87;
end 13'h14a7:    begin Red = 8'hd3;    Green = 8'had;    Blue = 8'h66;
end 13'h14a8:    begin Red = 8'hac;    Green = 8'h83;    Blue = 8'h57;
end 13'h14a9:    begin Red = 8'hf3;    Green = 8'hc7;    Blue = 8'h8a;
end 13'h14aa:    begin Red = 8'heb;    Green = 8'hbd;    Blue = 8'h7f;
end 13'h14ab:    begin Red = 8'hdd;    Green = 8'hb1;    Blue = 8'h72;
end 13'h14ac:    begin Red = 8'hde;    Green = 8'hb5;    Blue = 8'h7d;
end 13'h14ad:    begin Red = 8'hb2;    Green = 8'h8f;    Blue = 8'h59;
end 13'h14ae:    begin Red = 8'hd3;    Green = 8'hac;    Blue = 8'h71;
end 13'h14af:    begin Red = 8'hd3;    Green = 8'ha9;    Blue = 8'h6d;
end 13'h14b0:    begin Red = 8'hd4;    Green = 8'ha2;    Blue = 8'h65;
end 13'h14b1:    begin Red = 8'hbc;    Green = 8'h9d;    Blue = 8'h67;
end 13'h14b2:    begin Red = 8'ha2;    Green = 8'h7e;    Blue = 8'h4a;
end 13'h14b3:    begin Red = 8'haf;    Green = 8'h8f;    Blue = 8'h60;
end 13'h14b4:    begin Red = 8'hf2;    Green = 8'hec;    Blue = 8'hba;
end 13'h14b5:    begin Red = 8'hef;    Green = 8'hef;    Blue = 8'hb9;
end 13'h14b6:    begin Red = 8'hed;    Green = 8'he3;    Blue = 8'hb0;
end 13'h14b7:    begin Red = 8'hff;    Green = 8'hff;    Blue = 8'hd2;
end 13'h14b8:    begin Red = 8'hfb;    Green = 8'hff;    Blue = 8'hd5;
end 13'h14b9:    begin Red = 8'hfa;    Green = 8'hfd;    Blue = 8'hd0;
end 13'h14ba:    begin Red = 8'hfa;    Green = 8'hfe;    Blue = 8'hcb;
end 13'h14bb:    begin Red = 8'hfe;    Green = 8'hfc;    Blue = 8'hd5;
end 13'h14bc:    begin Red = 8'he4;    Green = 8'hd9;    Blue = 8'hab;
end 13'h14bd:    begin Red = 8'hfd;    Green = 8'hff;    Blue = 8'hce;
end 13'h14be:    begin Red = 8'hf8;    Green = 8'hff;    Blue = 8'hd2;
end 13'h14bf:    begin Red = 8'hf7;    Green = 8'heb;    Blue = 8'hc3;
end 13'h14c0:    begin Red = 8'hed;    Green = 8'he8;    Blue = 8'hae;
end 13'h14c1:    begin Red = 8'he8;    Green = 8'he7;    Blue = 8'hb9;
end 13'h14c2:    begin Red = 8'h98;    Green = 8'ha7;    Blue = 8'h8f;
end 13'h14c3:    begin Red = 8'h52;    Green = 8'h53;    Blue = 8'h55;
end 13'h14c4:    begin Red = 8'h64;    Green = 8'h68;    Blue = 8'h67;
end 13'h14c5:    begin Red = 8'h78;    Green = 8'h6c;    Blue = 8'h6e;
end 13'h14c6:    begin Red = 8'h00;    Green = 8'h04;    Blue = 8'h00;
end 13'h14c7:    begin Red = 8'h96;    Green = 8'h73;    Blue = 8'h9a;
end 13'h14c8:    begin Red = 8'h98;    Green = 8'h6e;    Blue = 8'h8c;
end 13'h14c9:    begin Red = 8'hb6;    Green = 8'h7f;    Blue = 8'hab;
end 13'h14ca:    begin Red = 8'hd7;    Green = 8'hb8;    Blue = 8'h65;
end 13'h14cb:    begin Red = 8'ha8;    Green = 8'h8a;    Blue = 8'h50;
end 13'h14cc:    begin Red = 8'h84;    Green = 8'h81;    Blue = 8'h7a;
end 13'h14cd:    begin Red = 8'h8a;    Green = 8'h87;    Blue = 8'h80;
end 13'h14ce:    begin Red = 8'heb;    Green = 8'hc3;    Blue = 8'h85;
end 13'h14cf:    begin Red = 8'hd9;    Green = 8'hae;    Blue = 8'h69;
end 13'h14d0:    begin Red = 8'hc2;    Green = 8'h99;    Blue = 8'h65;
end 13'h14d1:    begin Red = 8'h40;    Green = 8'h2e;    Blue = 8'h24;
end 13'h14d2:    begin Red = 8'h4e;    Green = 8'h3b;    Blue = 8'h2d;
end 13'h14d3:    begin Red = 8'h78;    Green = 8'h62;    Blue = 8'h4a;
end 13'h14d4:    begin Red = 8'h76;    Green = 8'h5e;    Blue = 8'h46;
end 13'h14d5:    begin Red = 8'h75;    Green = 8'h5d;    Blue = 8'h41;
end 13'h14d6:    begin Red = 8'hd8;    Green = 8'hb1;    Blue = 8'h64;
end 13'h14d7:    begin Red = 8'he3;    Green = 8'hb6;    Blue = 8'h7b;
end 13'h14d8:    begin Red = 8'h4e;    Green = 8'h33;    Blue = 8'h2a;
end 13'h14d9:    begin Red = 8'h46;    Green = 8'h32;    Blue = 8'h27;
end 13'h14da:    begin Red = 8'h43;    Green = 8'h2b;    Blue = 8'h1e;
end 13'h14db:    begin Red = 8'h69;    Green = 8'h53;    Blue = 8'h3c;
end 13'h14dc:    begin Red = 8'h64;    Green = 8'h4e;    Blue = 8'h39;
end 13'h14dd:    begin Red = 8'hdd;    Green = 8'hea;    Blue = 8'hca;
end 13'h14de:    begin Red = 8'hdd;    Green = 8'hdf;    Blue = 8'hbd;
end 13'h14df:    begin Red = 8'h9a;    Green = 8'ha5;    Blue = 8'h90;
end 13'h14e0:    begin Red = 8'h9f;    Green = 8'ha8;    Blue = 8'h97;
end 13'h14e1:    begin Red = 8'h5d;    Green = 8'h4b;    Blue = 8'h35;
end 13'h14e2:    begin Red = 8'h57;    Green = 8'h46;    Blue = 8'h34;
end 13'h14e3:    begin Red = 8'hb2;    Green = 8'h92;    Blue = 8'h61;
end 13'h14e4:    begin Red = 8'hce;    Green = 8'hc5;    Blue = 8'h9c;
end 13'h14e5:    begin Red = 8'heb;    Green = 8'he1;    Blue = 8'hbd;
end 13'h14e6:    begin Red = 8'h63;    Green = 8'h5f;    Blue = 8'h5e;
end 13'h14e7:    begin Red = 8'h83;    Green = 8'h79;    Blue = 8'h77;
end 13'h14e8:    begin Red = 8'h24;    Green = 8'h1e;    Blue = 8'h12;
end 13'h14e9:    begin Red = 8'h99;    Green = 8'h7c;    Blue = 8'h96;
end 13'h14ea:    begin Red = 8'h9a;    Green = 8'h75;    Blue = 8'h8e;
end 13'h14eb:    begin Red = 8'haf;    Green = 8'h84;    Blue = 8'ha6;
end 13'h14ec:    begin Red = 8'had;    Green = 8'hb3;    Blue = 8'h9a;
end 13'h14ed:    begin Red = 8'h3e;    Green = 8'h36;    Blue = 8'h36;
end 13'h14ee:    begin Red = 8'hd2;    Green = 8'hb3;    Blue = 8'h66;
end 13'h14ef:    begin Red = 8'hc5;    Green = 8'haa;    Blue = 8'h6f;
end 13'h14f0:    begin Red = 8'h82;    Green = 8'h7f;    Blue = 8'h7e;
end 13'h14f1:    begin Red = 8'h41;    Green = 8'h37;    Blue = 8'h3a;
end 13'h14f2:    begin Red = 8'h3f;    Green = 8'h38;    Blue = 8'h34;
end 13'h14f3:    begin Red = 8'hd4;    Green = 8'ha4;    Blue = 8'h62;
end 13'h14f4:    begin Red = 8'he8;    Green = 8'hbb;    Blue = 8'h7a;
end 13'h14f5:    begin Red = 8'hd9;    Green = 8'ha7;    Blue = 8'h6a;
end 13'h14f6:    begin Red = 8'h4d;    Green = 8'h30;    Blue = 8'h1e;
end 13'h14f7:    begin Red = 8'h5d;    Green = 8'h44;    Blue = 8'h2e;
end 13'h14f8:    begin Red = 8'h90;    Green = 8'h74;    Blue = 8'h4d;
end 13'h14f9:    begin Red = 8'h86;    Green = 8'h6a;    Blue = 8'h45;
end 13'h14fa:    begin Red = 8'h87;    Green = 8'h6f;    Blue = 8'h4d;
end 13'h14fb:    begin Red = 8'h85;    Green = 8'h6b;    Blue = 8'h48;
end 13'h14fc:    begin Red = 8'h83;    Green = 8'h69;    Blue = 8'h46;
end 13'h14fd:    begin Red = 8'hcf;    Green = 8'h9f;    Blue = 8'h61;
end 13'h14fe:    begin Red = 8'he6;    Green = 8'hb8;    Blue = 8'h7c;
end 13'h14ff:    begin Red = 8'he0;    Green = 8'hb7;    Blue = 8'h77;
end 13'h1500:    begin Red = 8'hca;    Green = 8'h9e;    Blue = 8'h5d;
end 13'h1501:    begin Red = 8'h50;    Green = 8'h3b;    Blue = 8'h26;
end 13'h1502:    begin Red = 8'h7e;    Green = 8'h6b;    Blue = 8'h43;
end 13'h1503:    begin Red = 8'h77;    Green = 8'h60;    Blue = 8'h41;
end 13'h1504:    begin Red = 8'h79;    Green = 8'h62;    Blue = 8'h43;
end 13'h1505:    begin Red = 8'h73;    Green = 8'h5a;    Blue = 8'h3c;
end 13'h1506:    begin Red = 8'hdd;    Green = 8'he7;    Blue = 8'hc5;
end 13'h1507:    begin Red = 8'h73;    Green = 8'h59;    Blue = 8'h40;
end 13'h1508:    begin Red = 8'h6f;    Green = 8'h5c;    Blue = 8'h3b;
end 13'h1509:    begin Red = 8'h6a;    Green = 8'h56;    Blue = 8'h3b;
end 13'h150a:    begin Red = 8'ha6;    Green = 8'h8b;    Blue = 8'h60;
end 13'h150b:    begin Red = 8'hfd;    Green = 8'he8;    Blue = 8'hbb;
end 13'h150c:    begin Red = 8'hbd;    Green = 8'h9d;    Blue = 8'h74;
end 13'h150d:    begin Red = 8'hb7;    Green = 8'h8e;    Blue = 8'h60;
end 13'h150e:    begin Red = 8'h27;    Green = 8'h20;    Blue = 8'h18;
end 13'h150f:    begin Red = 8'h32;    Green = 8'h28;    Blue = 8'h1f;
end 13'h1510:    begin Red = 8'h9a;    Green = 8'h76;    Blue = 8'h95;
end 13'h1511:    begin Red = 8'h9b;    Green = 8'h6d;    Blue = 8'h99;
end 13'h1512:    begin Red = 8'hc9;    Green = 8'ha6;    Blue = 8'h5f;
end 13'h1513:    begin Red = 8'hb7;    Green = 8'h9d;    Blue = 8'h5b;
end 13'h1514:    begin Red = 8'hc7;    Green = 8'hab;    Blue = 8'h5e;
end 13'h1515:    begin Red = 8'hcf;    Green = 8'haf;    Blue = 8'h6f;
end 13'h1516:    begin Red = 8'h80;    Green = 8'h78;    Blue = 8'h68;
end 13'h1517:    begin Red = 8'heb;    Green = 8'he6;    Blue = 8'hcd;
end 13'h1518:    begin Red = 8'he0;    Green = 8'hbd;    Blue = 8'h87;
end 13'h1519:    begin Red = 8'hf4;    Green = 8'hd1;    Blue = 8'h9b;
end 13'h151a:    begin Red = 8'hf0;    Green = 8'hcf;    Blue = 8'h9a;
end 13'h151b:    begin Red = 8'hcd;    Green = 8'hb0;    Blue = 8'h78;
end 13'h151c:    begin Red = 8'h62;    Green = 8'h48;    Blue = 8'h31;
end 13'h151d:    begin Red = 8'h8b;    Green = 8'h71;    Blue = 8'h4e;
end 13'h151e:    begin Red = 8'h9a;    Green = 8'h80;    Blue = 8'h5d;
end 13'h151f:    begin Red = 8'h9c;    Green = 8'h82;    Blue = 8'h5f;
end 13'h1520:    begin Red = 8'h87;    Green = 8'h68;    Blue = 8'h49;
end 13'h1521:    begin Red = 8'hf3;    Green = 8'hcd;    Blue = 8'h8e;
end 13'h1522:    begin Red = 8'hdb;    Green = 8'hba;    Blue = 8'h85;
end 13'h1523:    begin Red = 8'he1;    Green = 8'hc6;    Blue = 8'h8f;
end 13'h1524:    begin Red = 8'h83;    Green = 8'h68;    Blue = 8'h4d;
end 13'h1525:    begin Red = 8'h81;    Green = 8'h6c;    Blue = 8'h4f;
end 13'h1526:    begin Red = 8'h79;    Green = 8'h65;    Blue = 8'h4d;
end 13'h1527:    begin Red = 8'hb9;    Green = 8'h9d;    Blue = 8'h75;
end 13'h1528:    begin Red = 8'hb6;    Green = 8'h9f;    Blue = 8'h75;
end 13'h1529:    begin Red = 8'ha0;    Green = 8'h93;    Blue = 8'h4f;
end 13'h152a:    begin Red = 8'ha4;    Green = 8'h87;    Blue = 8'h4b;
end 13'h152b:    begin Red = 8'ha3;    Green = 8'h8e;    Blue = 8'h4d;
end 13'h152c:    begin Red = 8'hc3;    Green = 8'ha8;    Blue = 8'h63;
end 13'h152d:    begin Red = 8'hbc;    Green = 8'ha4;    Blue = 8'h5a;
end 13'h152e:    begin Red = 8'hc8;    Green = 8'hab;    Blue = 8'h65;
end 13'h152f:    begin Red = 8'hc6;    Green = 8'hb0;    Blue = 8'h67;
end 13'h1530:    begin Red = 8'hde;    Green = 8'hda;    Blue = 8'haa;
end 13'h1531:    begin Red = 8'hd1;    Green = 8'hd4;    Blue = 8'ha9;
end 13'h1532:    begin Red = 8'hfb;    Green = 8'hfd;    Blue = 8'hd8;
end 13'h1533:    begin Red = 8'hfc;    Green = 8'hfd;    Blue = 8'hd3;
end 13'h1534:    begin Red = 8'hfe;    Green = 8'hec;    Blue = 8'hba;
end 13'h1535:    begin Red = 8'ha1;    Green = 8'h88;    Blue = 8'h45;
end 13'h1536:    begin Red = 8'h9f;    Green = 8'h8c;    Blue = 8'h48;
end 13'h1537:    begin Red = 8'ha0;    Green = 8'h88;    Blue = 8'h4a;
end 13'h1538:    begin Red = 8'hd4;    Green = 8'he4;    Blue = 8'hbd;
end 13'h1539:    begin Red = 8'hb7;    Green = 8'ha3;    Blue = 8'h5c;
end 13'h153a:    begin Red = 8'hbe;    Green = 8'ha6;    Blue = 8'h60;
end 13'h153b:    begin Red = 8'hbd;    Green = 8'had;    Blue = 8'h62;
end 13'h153c:    begin Red = 8'hb9;    Green = 8'ha3;    Blue = 8'h58;
end 13'h153d:    begin Red = 8'hc0;    Green = 8'ha9;    Blue = 8'h59;
end 13'h153e:    begin Red = 8'hc9;    Green = 8'hb1;    Blue = 8'h6b;
end 13'h153f:    begin Red = 8'hc7;    Green = 8'ha9;    Blue = 8'h63;
end 13'h1540:    begin Red = 8'hcb;    Green = 8'haf;    Blue = 8'h66;
end 13'h1541:    begin Red = 8'hb9;    Green = 8'h95;    Blue = 8'h49;
end 13'h1542:    begin Red = 8'h24;    Green = 8'h24;    Blue = 8'h18;
end 13'h1543:    begin Red = 8'h32;    Green = 8'h25;    Blue = 8'h1c;
end 13'h1544:    begin Red = 8'haf;    Green = 8'h88;    Blue = 8'ha5;
end 13'h1545:    begin Red = 8'h98;    Green = 8'h78;    Blue = 8'h90;
end 13'h1546:    begin Red = 8'hb2;    Green = 8'ha6;    Blue = 8'ha3;
end 13'h1547:    begin Red = 8'hff;    Green = 8'hfa;    Blue = 8'he4;
end 13'h1548:    begin Red = 8'hff;    Green = 8'hf6;    Blue = 8'he2;
end 13'h1549:    begin Red = 8'hc4;    Green = 8'ha7;    Blue = 8'h67;
end 13'h154a:    begin Red = 8'h72;    Green = 8'h69;    Blue = 8'h65;
end 13'h154b:    begin Red = 8'hbb;    Green = 8'h9d;    Blue = 8'h61;
end 13'h154c:    begin Red = 8'h92;    Green = 8'h84;    Blue = 8'h74;
end 13'h154d:    begin Red = 8'hbf;    Green = 8'hc7;    Blue = 8'hc7;
end 13'h154e:    begin Red = 8'he5;    Green = 8'hf0;    Blue = 8'he2;
end 13'h154f:    begin Red = 8'hf6;    Green = 8'hd5;    Blue = 8'ha2;
end 13'h1550:    begin Red = 8'hf1;    Green = 8'hd0;    Blue = 8'h9d;
end 13'h1551:    begin Red = 8'hf6;    Green = 8'hd0;    Blue = 8'h9f;
end 13'h1552:    begin Red = 8'he3;    Green = 8'hc5;    Blue = 8'h91;
end 13'h1553:    begin Red = 8'h50;    Green = 8'h4d;    Blue = 8'h3e;
end 13'h1554:    begin Red = 8'h9f;    Green = 8'h85;    Blue = 8'h62;
end 13'h1555:    begin Red = 8'hf6;    Green = 8'hca;    Blue = 8'h8b;
end 13'h1556:    begin Red = 8'h5a;    Green = 8'h40;    Blue = 8'h2f;
end 13'h1557:    begin Red = 8'h97;    Green = 8'h7c;    Blue = 8'h61;
end 13'h1558:    begin Red = 8'h8f;    Green = 8'h70;    Blue = 8'h54;
end 13'h1559:    begin Red = 8'h87;    Green = 8'h70;    Blue = 8'h51;
end 13'h155a:    begin Red = 8'he2;    Green = 8'hec;    Blue = 8'hca;
end 13'h155b:    begin Red = 8'hc2;    Green = 8'h9e;    Blue = 8'h6c;
end 13'h155c:    begin Red = 8'hb0;    Green = 8'h99;    Blue = 8'h6d;
end 13'h155d:    begin Red = 8'hbf;    Green = 8'ha7;    Blue = 8'h7b;
end 13'h155e:    begin Red = 8'hc1;    Green = 8'ha3;    Blue = 8'h7f;
end 13'h155f:    begin Red = 8'h9a;    Green = 8'h7f;    Blue = 8'h61;
end 13'h1560:    begin Red = 8'hc2;    Green = 8'h87;    Blue = 8'hb3;
end 13'h1561:    begin Red = 8'hc9;    Green = 8'h8c;    Blue = 8'hb6;
end 13'h1562:    begin Red = 8'h9e;    Green = 8'h74;    Blue = 8'h98;
end 13'h1563:    begin Red = 8'ha6;    Green = 8'h78;    Blue = 8'h9c;
end 13'h1564:    begin Red = 8'hbf;    Green = 8'h84;    Blue = 8'hb4;
end 13'h1565:    begin Red = 8'ha4;    Green = 8'h72;    Blue = 8'h97;
end 13'h1566:    begin Red = 8'ha8;    Green = 8'h74;    Blue = 8'h98;
end 13'h1567:    begin Red = 8'ha2;    Green = 8'h74;    Blue = 8'h99;
end 13'h1568:    begin Red = 8'h94;    Green = 8'h64;    Blue = 8'h8a;
end 13'h1569:    begin Red = 8'h97;    Green = 8'h67;    Blue = 8'h8f;
end 13'h156a:    begin Red = 8'h78;    Green = 8'h53;    Blue = 8'h75;
end 13'h156b:    begin Red = 8'h84;    Green = 8'h58;    Blue = 8'h79;
end 13'h156c:    begin Red = 8'h7d;    Green = 8'h50;    Blue = 8'h77;
end 13'h156d:    begin Red = 8'h9e;    Green = 8'h68;    Blue = 8'h88;
end 13'h156e:    begin Red = 8'hbf;    Green = 8'h82;    Blue = 8'hbd;
end 13'h156f:    begin Red = 8'hc4;    Green = 8'h85;    Blue = 8'hba;
end 13'h1570:    begin Red = 8'hc1;    Green = 8'h86;    Blue = 8'hbc;
end 13'h1571:    begin Red = 8'h9d;    Green = 8'h71;    Blue = 8'h95;
end 13'h1572:    begin Red = 8'h97;    Green = 8'h6e;    Blue = 8'h96;
end 13'h1573:    begin Red = 8'hc2;    Green = 8'h88;    Blue = 8'hb8;
end 13'h1574:    begin Red = 8'hc1;    Green = 8'h83;    Blue = 8'hb2;
end 13'h1575:    begin Red = 8'h92;    Green = 8'h60;    Blue = 8'h85;
end 13'h1576:    begin Red = 8'h96;    Green = 8'h66;    Blue = 8'h8c;
end 13'h1577:    begin Red = 8'h80;    Green = 8'h54;    Blue = 8'h75;
end 13'h1578:    begin Red = 8'h9d;    Green = 8'h69;    Blue = 8'h8f;
end 13'h1579:    begin Red = 8'h9c;    Green = 8'h65;    Blue = 8'h8f;
end 13'h157a:    begin Red = 8'ha1;    Green = 8'h6d;    Blue = 8'h93;
end 13'h157b:    begin Red = 8'h86;    Green = 8'h5a;    Blue = 8'h7b;
end 13'h157c:    begin Red = 8'h7f;    Green = 8'h55;    Blue = 8'h79;
end 13'h157d:    begin Red = 8'h9e;    Green = 8'h67;    Blue = 8'h91;
end 13'h157e:    begin Red = 8'h7e;    Green = 8'h59;    Blue = 8'h7a;
end 13'h157f:    begin Red = 8'h8c;    Green = 8'h50;    Blue = 8'h90;
end 13'h1580:    begin Red = 8'h38;    Green = 8'h30;    Blue = 8'h23;
end 13'h1581:    begin Red = 8'hf6;    Green = 8'hdb;    Blue = 8'hb0;
end 13'h1582:    begin Red = 8'h9b;    Green = 8'h78;    Blue = 8'h8a;
end 13'h1583:    begin Red = 8'h9e;    Green = 8'h79;    Blue = 8'h8e;
end 13'h1584:    begin Red = 8'hae;    Green = 8'h89;    Blue = 8'ha0;
end 13'h1585:    begin Red = 8'hac;    Green = 8'h95;    Blue = 8'h87;
end 13'h1586:    begin Red = 8'ha5;    Green = 8'h8c;    Blue = 8'h51;
end 13'h1587:    begin Red = 8'hea;    Green = 8'hde;    Blue = 8'hc5;
end 13'h1588:    begin Red = 8'h66;    Green = 8'h5d;    Blue = 8'h53;
end 13'h1589:    begin Red = 8'hf0;    Green = 8'hd8;    Blue = 8'hc5;
end 13'h158a:    begin Red = 8'hc2;    Green = 8'hc2;    Blue = 8'ha7;
end 13'h158b:    begin Red = 8'hd8;    Green = 8'h91;    Blue = 8'h34;
end 13'h158c:    begin Red = 8'hd7;    Green = 8'h95;    Blue = 8'h44;
end 13'h158d:    begin Red = 8'hd5;    Green = 8'h94;    Blue = 8'h41;
end 13'h158e:    begin Red = 8'hce;    Green = 8'h8e;    Blue = 8'h34;
end 13'h158f:    begin Red = 8'he6;    Green = 8'hc2;    Blue = 8'h86;
end 13'h1590:    begin Red = 8'h82;    Green = 8'h6e;    Blue = 8'h4b;
end 13'h1591:    begin Red = 8'hde;    Green = 8'had;    Blue = 8'h6a;
end 13'h1592:    begin Red = 8'he2;    Green = 8'hc4;    Blue = 8'h84;
end 13'h1593:    begin Red = 8'he1;    Green = 8'hba;    Blue = 8'h7f;
end 13'h1594:    begin Red = 8'hdd;    Green = 8'hb3;    Blue = 8'h77;
end 13'h1595:    begin Red = 8'hc6;    Green = 8'hd2;    Blue = 8'haf;
end 13'h1596:    begin Red = 8'hb2;    Green = 8'h8a;    Blue = 8'h56;
end 13'h1597:    begin Red = 8'h8f;    Green = 8'h69;    Blue = 8'h42;
end 13'h1598:    begin Red = 8'h7c;    Green = 8'h57;    Blue = 8'h79;
end 13'h1599:    begin Red = 8'h82;    Green = 8'h5a;    Blue = 8'h7c;
end 13'h159a:    begin Red = 8'h7f;    Green = 8'h58;    Blue = 8'h77;
end 13'h159b:    begin Red = 8'h76;    Green = 8'h56;    Blue = 8'h23;
end 13'h159c:    begin Red = 8'h85;    Green = 8'h6f;    Blue = 8'h3e;
end 13'h159d:    begin Red = 8'haf;    Green = 8'h82;    Blue = 8'h47;
end 13'h159e:    begin Red = 8'ha5;    Green = 8'h85;    Blue = 8'h48;
end 13'h159f:    begin Red = 8'ha1;    Green = 8'h83;    Blue = 8'h47;
end 13'h15a0:    begin Red = 8'ha6;    Green = 8'h83;    Blue = 8'h4b;
end 13'h15a1:    begin Red = 8'hae;    Green = 8'h7f;    Blue = 8'h51;
end 13'h15a2:    begin Red = 8'hfa;    Green = 8'he7;    Blue = 8'ha3;
end 13'h15a3:    begin Red = 8'h8e;    Green = 8'h61;    Blue = 8'h82;
end 13'h15a4:    begin Red = 8'h99;    Green = 8'h6b;    Blue = 8'h92;
end 13'h15a5:    begin Red = 8'h9e;    Green = 8'h6c;    Blue = 8'h92;
end 13'h15a6:    begin Red = 8'h85;    Green = 8'h4d;    Blue = 8'h8a;
end 13'h15a7:    begin Red = 8'h33;    Green = 8'h31;    Blue = 8'h22;
end 13'h15a8:    begin Red = 8'ha5;    Green = 8'h8d;    Blue = 8'h5d;
end 13'h15a9:    begin Red = 8'hd3;    Green = 8'hb3;    Blue = 8'h6d;
end 13'h15aa:    begin Red = 8'hcd;    Green = 8'hc6;    Blue = 8'had;
end 13'h15ab:    begin Red = 8'h94;    Green = 8'h84;    Blue = 8'h5c;
end 13'h15ac:    begin Red = 8'hb7;    Green = 8'hba;    Blue = 8'h98;
end 13'h15ad:    begin Red = 8'hf6;    Green = 8'hac;    Blue = 8'h42;
end 13'h15ae:    begin Red = 8'hcc;    Green = 8'h90;    Blue = 8'h3f;
end 13'h15af:    begin Red = 8'hd2;    Green = 8'h8c;    Blue = 8'h36;
end 13'h15b0:    begin Red = 8'h9b;    Green = 8'h7f;    Blue = 8'h5a;
end 13'h15b1:    begin Red = 8'h85;    Green = 8'h6f;    Blue = 8'h4a;
end 13'h15b2:    begin Red = 8'he5;    Green = 8'hb2;    Blue = 8'h71;
end 13'h15b3:    begin Red = 8'hdf;    Green = 8'hb5;    Blue = 8'h79;
end 13'h15b4:    begin Red = 8'hcd;    Green = 8'ha0;    Blue = 8'h65;
end 13'h15b5:    begin Red = 8'h87;    Green = 8'h5f;    Blue = 8'h82;
end 13'h15b6:    begin Red = 8'h85;    Green = 8'h5d;    Blue = 8'h80;
end 13'h15b7:    begin Red = 8'h8a;    Green = 8'h5c;    Blue = 8'h80;
end 13'h15b8:    begin Red = 8'ha8;    Green = 8'h6f;    Blue = 8'h98;
end 13'h15b9:    begin Red = 8'h9e;    Green = 8'h6e;    Blue = 8'h98;
end 13'h15ba:    begin Red = 8'ha7;    Green = 8'h75;    Blue = 8'h9b;
end 13'h15bb:    begin Red = 8'h7b;    Green = 8'h6f;    Blue = 8'h3f;
end 13'h15bc:    begin Red = 8'h9b;    Green = 8'h8a;    Blue = 8'h3c;
end 13'h15bd:    begin Red = 8'ha6;    Green = 8'h88;    Blue = 8'h3f;
end 13'h15be:    begin Red = 8'hb7;    Green = 8'h8f;    Blue = 8'h47;
end 13'h15bf:    begin Red = 8'hba;    Green = 8'h8a;    Blue = 8'h4a;
end 13'h15c0:    begin Red = 8'ha8;    Green = 8'h8e;    Blue = 8'h37;
end 13'h15c1:    begin Red = 8'ha8;    Green = 8'h8f;    Blue = 8'h3b;
end 13'h15c2:    begin Red = 8'hb1;    Green = 8'h8f;    Blue = 8'h47;
end 13'h15c3:    begin Red = 8'hbc;    Green = 8'h87;    Blue = 8'h43;
end 13'h15c4:    begin Red = 8'hac;    Green = 8'h8b;    Blue = 8'h44;
end 13'h15c5:    begin Red = 8'hb3;    Green = 8'h91;    Blue = 8'h49;
end 13'h15c6:    begin Red = 8'ha9;    Green = 8'h8a;    Blue = 8'h3a;
end 13'h15c7:    begin Red = 8'hae;    Green = 8'h87;    Blue = 8'h44;
end 13'h15c8:    begin Red = 8'hfc;    Green = 8'hec;    Blue = 8'hb0;
end 13'h15c9:    begin Red = 8'hc7;    Green = 8'h92;    Blue = 8'hc0;
end 13'h15ca:    begin Red = 8'h9b;    Green = 8'h6b;    Blue = 8'h95;
end 13'h15cb:    begin Red = 8'ha5;    Green = 8'h6d;    Blue = 8'h9a;
end 13'h15cc:    begin Red = 8'h82;    Green = 8'h5d;    Blue = 8'h7e;
end 13'h15cd:    begin Red = 8'ha5;    Green = 8'h6e;    Blue = 8'h96;
end 13'h15ce:    begin Red = 8'h8c;    Green = 8'h5e;    Blue = 8'h82;
end 13'h15cf:    begin Red = 8'h8d;    Green = 8'h53;    Blue = 8'h8e;
end 13'h15d0:    begin Red = 8'ha8;    Green = 8'h80;    Blue = 8'h9c;
end 13'h15d1:    begin Red = 8'haf;    Green = 8'hae;    Blue = 8'h9d;
end 13'h15d2:    begin Red = 8'hcf;    Green = 8'hb7;    Blue = 8'ha3;
end 13'h15d3:    begin Red = 8'h94;    Green = 8'h89;    Blue = 8'h59;
end 13'h15d4:    begin Red = 8'hd7;    Green = 8'hbc;    Blue = 8'h9f;
end 13'h15d5:    begin Red = 8'hbe;    Green = 8'hac;    Blue = 8'h84;
end 13'h15d6:    begin Red = 8'hb7;    Green = 8'ha6;    Blue = 8'h7e;
end 13'h15d7:    begin Red = 8'he0;    Green = 8'he4;    Blue = 8'hd4;
end 13'h15d8:    begin Red = 8'h5d;    Green = 8'h4d;    Blue = 8'h3e;
end 13'h15d9:    begin Red = 8'h82;    Green = 8'h6c;    Blue = 8'h47;
end 13'h15da:    begin Red = 8'he1;    Green = 8'hae;    Blue = 8'h6d;
end 13'h15db:    begin Red = 8'h59;    Green = 8'h40;    Blue = 8'h2a;
end 13'h15dc:    begin Red = 8'h7e;    Green = 8'h67;    Blue = 8'h48;
end 13'h15dd:    begin Red = 8'h77;    Green = 8'h4b;    Blue = 8'h6c;
end 13'h15de:    begin Red = 8'h81;    Green = 8'h4d;    Blue = 8'h74;
end 13'h15df:    begin Red = 8'h69;    Green = 8'h3d;    Blue = 8'h5e;
end 13'h15e0:    begin Red = 8'h64;    Green = 8'h3f;    Blue = 8'h60;
end 13'h15e1:    begin Red = 8'h61;    Green = 8'h3c;    Blue = 8'h5d;
end 13'h15e2:    begin Red = 8'h79;    Green = 8'h49;    Blue = 8'h6f;
end 13'h15e3:    begin Red = 8'h6a;    Green = 8'h41;    Blue = 8'h63;
end 13'h15e4:    begin Red = 8'h81;    Green = 8'h4a;    Blue = 8'h72;
end 13'h15e5:    begin Red = 8'h62;    Green = 8'h3b;    Blue = 8'h5a;
end 13'h15e6:    begin Red = 8'h61;    Green = 8'h3a;    Blue = 8'h57;
end 13'h15e7:    begin Red = 8'h94;    Green = 8'h69;    Blue = 8'h97;
end 13'h15e8:    begin Red = 8'hb0;    Green = 8'h6a;    Blue = 8'ha0;
end 13'h15e9:    begin Red = 8'h57;    Green = 8'h57;    Blue = 8'h59;
end 13'h15ea:    begin Red = 8'h55;    Green = 8'h5a;    Blue = 8'h54;
end 13'h15eb:    begin Red = 8'h99;    Green = 8'h68;    Blue = 8'h95;
end 13'h15ec:    begin Red = 8'h9e;    Green = 8'h64;    Blue = 8'h8c;
end 13'h15ed:    begin Red = 8'h58;    Green = 8'h57;    Blue = 8'h53;
end 13'h15ee:    begin Red = 8'h48;    Green = 8'h53;    Blue = 8'h4f;
end 13'h15ef:    begin Red = 8'ha2;    Green = 8'h66;    Blue = 8'h99;
end 13'h15f0:    begin Red = 8'h4d;    Green = 8'h52;    Blue = 8'h4c;
end 13'h15f1:    begin Red = 8'ha7;    Green = 8'h69;    Blue = 8'h9c;
end 13'h15f2:    begin Red = 8'h95;    Green = 8'h6a;    Blue = 8'h88;
end 13'h15f3:    begin Red = 8'hff;    Green = 8'hf7;    Blue = 8'hb9;
end 13'h15f4:    begin Red = 8'h7b;    Green = 8'h4b;    Blue = 8'h73;
end 13'h15f5:    begin Red = 8'h77;    Green = 8'h47;    Blue = 8'h6d;
end 13'h15f6:    begin Red = 8'h6a;    Green = 8'h3e;    Blue = 8'h61;
end 13'h15f7:    begin Red = 8'h7e;    Green = 8'h4f;    Blue = 8'h73;
end 13'h15f8:    begin Red = 8'h7d;    Green = 8'h48;    Blue = 8'h72;
end 13'h15f9:    begin Red = 8'h61;    Green = 8'h2b;    Blue = 8'h65;
end 13'h15fa:    begin Red = 8'h2f;    Green = 8'h24;    Blue = 8'h1e;
end 13'h15fb:    begin Red = 8'hcf;    Green = 8'haf;    Blue = 8'h76;
end 13'h15fc:    begin Red = 8'ha3;    Green = 8'ha7;    Blue = 8'h43;
end 13'h15fd:    begin Red = 8'hb0;    Green = 8'hbb;    Blue = 8'h67;
end 13'h15fe:    begin Red = 8'h99;    Green = 8'h88;    Blue = 8'h56;
end 13'h15ff:    begin Red = 8'h75;    Green = 8'h72;    Blue = 8'h56;
end 13'h1600:    begin Red = 8'hd3;    Green = 8'hcc;    Blue = 8'had;
end 13'h1601:    begin Red = 8'hb8;    Green = 8'hb3;    Blue = 8'h9e;
end 13'h1602:    begin Red = 8'hf6;    Green = 8'ha4;    Blue = 8'h34;
end 13'h1603:    begin Red = 8'h48;    Green = 8'h36;    Blue = 8'h28;
end 13'h1604:    begin Red = 8'h6b;    Green = 8'h57;    Blue = 8'h3e;
end 13'h1605:    begin Red = 8'h89;    Green = 8'h79;    Blue = 8'h3e;
end 13'h1606:    begin Red = 8'h84;    Green = 8'h78;    Blue = 8'h3c;
end 13'h1607:    begin Red = 8'ha5;    Green = 8'h91;    Blue = 8'h52;
end 13'h1608:    begin Red = 8'ha2;    Green = 8'h8a;    Blue = 8'h4c;
end 13'h1609:    begin Red = 8'ha2;    Green = 8'h89;    Blue = 8'h50;
end 13'h160a:    begin Red = 8'ha7;    Green = 8'h8f;    Blue = 8'h51;
end 13'h160b:    begin Red = 8'h8c;    Green = 8'h6e;    Blue = 8'h3a;
end 13'h160c:    begin Red = 8'h49;    Green = 8'h56;    Blue = 8'h4c;
end 13'h160d:    begin Red = 8'h5e;    Green = 8'h55;    Blue = 8'h58;
end 13'h160e:    begin Red = 8'h49;    Green = 8'h4c;    Blue = 8'h41;
end 13'h160f:    begin Red = 8'h5a;    Green = 8'h57;    Blue = 8'h62;
end 13'h1610:    begin Red = 8'h42;    Green = 8'h50;    Blue = 8'h51;
end 13'h1611:    begin Red = 8'hab;    Green = 8'h6b;    Blue = 8'ha7;
end 13'h1612:    begin Red = 8'hb4;    Green = 8'h6c;    Blue = 8'h9e;
end 13'h1613:    begin Red = 8'h96;    Green = 8'h72;    Blue = 8'h38;
end 13'h1614:    begin Red = 8'h83;    Green = 8'h72;    Blue = 8'h3a;
end 13'h1615:    begin Red = 8'h86;    Green = 8'h76;    Blue = 8'h3a;
end 13'h1616:    begin Red = 8'h8b;    Green = 8'h7b;    Blue = 8'h3d;
end 13'h1617:    begin Red = 8'h9f;    Green = 8'h8b;    Blue = 8'h4e;
end 13'h1618:    begin Red = 8'ha2;    Green = 8'h8e;    Blue = 8'h51;
end 13'h1619:    begin Red = 8'ha6;    Green = 8'h89;    Blue = 8'h4d;
end 13'h161a:    begin Red = 8'h8c;    Green = 8'h73;    Blue = 8'h3d;
end 13'h161b:    begin Red = 8'h67;    Green = 8'h64;    Blue = 8'h51;
end 13'h161c:    begin Red = 8'h22;    Green = 8'h20;    Blue = 8'h14;
end 13'h161d:    begin Red = 8'hf3;    Green = 8'hdb;    Blue = 8'hab;
end 13'h161e:    begin Red = 8'h96;    Green = 8'h78;    Blue = 8'h93;
end 13'h161f:    begin Red = 8'h9b;    Green = 8'h7b;    Blue = 8'h90;
end 13'h1620:    begin Red = 8'ha0;    Green = 8'h84;    Blue = 8'h4b;
end 13'h1621:    begin Red = 8'hb2;    Green = 8'h97;    Blue = 8'h66;
end 13'h1622:    begin Red = 8'hb4;    Green = 8'h9b;    Blue = 8'h5c;
end 13'h1623:    begin Red = 8'h9c;    Green = 8'ha3;    Blue = 8'h34;
end 13'h1624:    begin Red = 8'h98;    Green = 8'h8c;    Blue = 8'h55;
end 13'h1625:    begin Red = 8'h9c;    Green = 8'h8d;    Blue = 8'h5e;
end 13'h1626:    begin Red = 8'h56;    Green = 8'h55;    Blue = 8'h34;
end 13'h1627:    begin Red = 8'hbb;    Green = 8'hc8;    Blue = 8'ha7;
end 13'h1628:    begin Red = 8'haf;    Green = 8'hb2;    Blue = 8'h8e;
end 13'h1629:    begin Red = 8'hfc;    Green = 8'ha3;    Blue = 8'h34;
end 13'h162a:    begin Red = 8'hf7;    Green = 8'ha9;    Blue = 8'h34;
end 13'h162b:    begin Red = 8'heb;    Green = 8'ha9;    Blue = 8'h40;
end 13'h162c:    begin Red = 8'hf3;    Green = 8'hae;    Blue = 8'h3f;
end 13'h162d:    begin Red = 8'hc9;    Green = 8'h8d;    Blue = 8'h3d;
end 13'h162e:    begin Red = 8'hd3;    Green = 8'h95;    Blue = 8'h3d;
end 13'h162f:    begin Red = 8'hce;    Green = 8'h94;    Blue = 8'h45;
end 13'h1630:    begin Red = 8'hcb;    Green = 8'h8d;    Blue = 8'h35;
end 13'h1631:    begin Red = 8'ha9;    Green = 8'h93;    Blue = 8'h5a;
end 13'h1632:    begin Red = 8'hdb;    Green = 8'hb3;    Blue = 8'h6e;
end 13'h1633:    begin Red = 8'hff;    Green = 8'hdb;    Blue = 8'h97;
end 13'h1634:    begin Red = 8'hfe;    Green = 8'hd1;    Blue = 8'h8d;
end 13'h1635:    begin Red = 8'hff;    Green = 8'hce;    Blue = 8'h8c;
end 13'h1636:    begin Red = 8'hfb;    Green = 8'hce;    Blue = 8'h8d;
end 13'h1637:    begin Red = 8'hd6;    Green = 8'ha1;    Blue = 8'h5b;
end 13'h1638:    begin Red = 8'hcb;    Green = 8'ha1;    Blue = 8'h59;
end 13'h1639:    begin Red = 8'ha8;    Green = 8'h8a;    Blue = 8'h56;
end 13'h163a:    begin Red = 8'hc9;    Green = 8'ha5;    Blue = 8'h67;
end 13'h163b:    begin Red = 8'hf0;    Green = 8'hc5;    Blue = 8'h80;
end 13'h163c:    begin Red = 8'he4;    Green = 8'hb8;    Blue = 8'h71;
end 13'h163d:    begin Red = 8'he5;    Green = 8'hb9;    Blue = 8'h78;
end 13'h163e:    begin Red = 8'hbb;    Green = 8'hc6;    Blue = 8'ha3;
end 13'h163f:    begin Red = 8'hb3;    Green = 8'hbe;    Blue = 8'h91;
end 13'h1640:    begin Red = 8'hde;    Green = 8'hac;    Blue = 8'h7b;
end 13'h1641:    begin Red = 8'hd0;    Green = 8'haa;    Blue = 8'h69;
end 13'h1642:    begin Red = 8'h86;    Green = 8'h6f;    Blue = 8'h46;
end 13'h1643:    begin Red = 8'h9b;    Green = 8'h80;    Blue = 8'h53;
end 13'h1644:    begin Red = 8'h97;    Green = 8'h7f;    Blue = 8'h53;
end 13'h1645:    begin Red = 8'h95;    Green = 8'h7d;    Blue = 8'h4f;
end 13'h1646:    begin Red = 8'h85;    Green = 8'h72;    Blue = 8'h37;
end 13'h1647:    begin Red = 8'h59;    Green = 8'h5c;    Blue = 8'h55;
end 13'h1648:    begin Red = 8'h42;    Green = 8'h59;    Blue = 8'h53;
end 13'h1649:    begin Red = 8'h5a;    Green = 8'h55;    Blue = 8'h52;
end 13'h164a:    begin Red = 8'h5a;    Green = 8'h59;    Blue = 8'h5e;
end 13'h164b:    begin Red = 8'h50;    Green = 8'h5d;    Blue = 8'h4c;
end 13'h164c:    begin Red = 8'h93;    Green = 8'h68;    Blue = 8'h93;
end 13'h164d:    begin Red = 8'h62;    Green = 8'h59;    Blue = 8'h54;
end 13'h164e:    begin Red = 8'ha1;    Green = 8'h6c;    Blue = 8'h9a;
end 13'h164f:    begin Red = 8'ha8;    Green = 8'h6d;    Blue = 8'h9d;
end 13'h1650:    begin Red = 8'h82;    Green = 8'h6c;    Blue = 8'h3d;
end 13'h1651:    begin Red = 8'h9d;    Green = 8'h7e;    Blue = 8'h52;
end 13'h1652:    begin Red = 8'h9c;    Green = 8'h81;    Blue = 8'h56;
end 13'h1653:    begin Red = 8'h9c;    Green = 8'h7b;    Blue = 8'h4e;
end 13'h1654:    begin Red = 8'h9a;    Green = 8'h7d;    Blue = 8'h45;
end 13'h1655:    begin Red = 8'h28;    Green = 8'h27;    Blue = 8'h15;
end 13'h1656:    begin Red = 8'hb2;    Green = 8'h86;    Blue = 8'ha5;
end 13'h1657:    begin Red = 8'ha1;    Green = 8'h7a;    Blue = 8'h91;
end 13'h1658:    begin Red = 8'had;    Green = 8'h85;    Blue = 8'ha1;
end 13'h1659:    begin Red = 8'h78;    Green = 8'h6e;    Blue = 8'h50;
end 13'h165a:    begin Red = 8'hbc;    Green = 8'ha7;    Blue = 8'h5e;
end 13'h165b:    begin Red = 8'h88;    Green = 8'h80;    Blue = 8'h78;
end 13'h165c:    begin Red = 8'hac;    Green = 8'hb2;    Blue = 8'h5a;
end 13'h165d:    begin Red = 8'h94;    Green = 8'h8b;    Blue = 8'h5e;
end 13'h165e:    begin Red = 8'hba;    Green = 8'hc9;    Blue = 8'h9d;
end 13'h165f:    begin Red = 8'hb1;    Green = 8'hb6;    Blue = 8'h9b;
end 13'h1660:    begin Red = 8'hf8;    Green = 8'hb0;    Blue = 8'h42;
end 13'h1661:    begin Red = 8'hf6;    Green = 8'hae;    Blue = 8'h46;
end 13'h1662:    begin Red = 8'hf9;    Green = 8'haa;    Blue = 8'h47;
end 13'h1663:    begin Red = 8'hca;    Green = 8'h94;    Blue = 8'h41;
end 13'h1664:    begin Red = 8'hcf;    Green = 8'h90;    Blue = 8'h46;
end 13'h1665:    begin Red = 8'hd9;    Green = 8'haa;    Blue = 8'h76;
end 13'h1666:    begin Red = 8'hd1;    Green = 8'hac;    Blue = 8'h75;
end 13'h1667:    begin Red = 8'hcc;    Green = 8'ha9;    Blue = 8'h73;
end 13'h1668:    begin Red = 8'hc6;    Green = 8'ha0;    Blue = 8'h61;
end 13'h1669:    begin Red = 8'hbf;    Green = 8'h9b;    Blue = 8'h6b;
end 13'h166a:    begin Red = 8'hb9;    Green = 8'ha0;    Blue = 8'h78;
end 13'h166b:    begin Red = 8'h88;    Green = 8'h6e;    Blue = 8'h3d;
end 13'h166c:    begin Red = 8'ha7;    Green = 8'h83;    Blue = 8'h47;
end 13'h166d:    begin Red = 8'hfd;    Green = 8'he0;    Blue = 8'hb4;
end 13'h166e:    begin Red = 8'h87;    Green = 8'h66;    Blue = 8'h80;
end 13'h166f:    begin Red = 8'h84;    Green = 8'h63;    Blue = 8'h7e;
end 13'h1670:    begin Red = 8'hac;    Green = 8'hb0;    Blue = 8'h61;
end 13'h1671:    begin Red = 8'h91;    Green = 8'h7f;    Blue = 8'h57;
end 13'h1672:    begin Red = 8'h95;    Green = 8'h88;    Blue = 8'h5f;
end 13'h1673:    begin Red = 8'h77;    Green = 8'h70;    Blue = 8'h57;
end 13'h1674:    begin Red = 8'hb4;    Green = 8'hbe;    Blue = 8'h9a;
end 13'h1675:    begin Red = 8'hf4;    Green = 8'hac;    Blue = 8'h3b;
end 13'h1676:    begin Red = 8'hfe;    Green = 8'hb9;    Blue = 8'h3c;
end 13'h1677:    begin Red = 8'hfe;    Green = 8'hb7;    Blue = 8'h36;
end 13'h1678:    begin Red = 8'hf4;    Green = 8'ha9;    Blue = 8'h46;
end 13'h1679:    begin Red = 8'he2;    Green = 8'h9e;    Blue = 8'h3a;
end 13'h167a:    begin Red = 8'hd2;    Green = 8'h99;    Blue = 8'h43;
end 13'h167b:    begin Red = 8'h75;    Green = 8'h61;    Blue = 8'h4b;
end 13'h167c:    begin Red = 8'h9b;    Green = 8'h75;    Blue = 8'h44;
end 13'h167d:    begin Red = 8'he2;    Green = 8'hb0;    Blue = 8'h73;
end 13'h167e:    begin Red = 8'h92;    Green = 8'h69;    Blue = 8'h3d;
end 13'h167f:    begin Red = 8'ha0;    Green = 8'h80;    Blue = 8'h4d;
end 13'h1680:    begin Red = 8'hc0;    Green = 8'h92;    Blue = 8'h5e;
end 13'h1681:    begin Red = 8'hbb;    Green = 8'h93;    Blue = 8'h58;
end 13'h1682:    begin Red = 8'hd8;    Green = 8'he2;    Blue = 8'hc3;
end 13'h1683:    begin Red = 8'hae;    Green = 8'h84;    Blue = 8'h52;
end 13'h1684:    begin Red = 8'ha5;    Green = 8'h80;    Blue = 8'h53;
end 13'h1685:    begin Red = 8'h00;    Green = 8'h01;    Blue = 8'h0b;
end 13'h1686:    begin Red = 8'h1c;    Green = 8'h18;    Blue = 8'h27;
end 13'h1687:    begin Red = 8'h01;    Green = 8'h3d;    Blue = 8'h19;
end 13'h1688:    begin Red = 8'h11;    Green = 8'h10;    Blue = 8'h18;
end 13'h1689:    begin Red = 8'h24;    Green = 8'h1e;    Blue = 8'h2c;
end 13'h168a:    begin Red = 8'h22;    Green = 8'h1f;    Blue = 8'h28;
end 13'h168b:    begin Red = 8'h25;    Green = 8'h1a;    Blue = 8'h2b;
end 13'h168c:    begin Red = 8'h00;    Green = 8'h10;    Blue = 8'h11;
end 13'h168d:    begin Red = 8'hed;    Green = 8'hd9;    Blue = 8'ha4;
end 13'h168e:    begin Red = 8'hec;    Green = 8'hda;    Blue = 8'hc8;
end 13'h168f:    begin Red = 8'hee;    Green = 8'hed;    Blue = 8'hd5;
end 13'h1690:    begin Red = 8'h95;    Green = 8'h65;    Blue = 8'h4a;
end 13'h1691:    begin Red = 8'h7f;    Green = 8'h6d;    Blue = 8'h3e;
end 13'h1692:    begin Red = 8'h9e;    Green = 8'h90;    Blue = 8'h5d;
end 13'h1693:    begin Red = 8'h69;    Green = 8'h64;    Blue = 8'h41;
end 13'h1694:    begin Red = 8'hbd;    Green = 8'hb7;    Blue = 8'h93;
end 13'h1695:    begin Red = 8'h98;    Green = 8'h81;    Blue = 8'h60;
end 13'h1696:    begin Red = 8'h8a;    Green = 8'h70;    Blue = 8'h54;
end 13'h1697:    begin Red = 8'hc1;    Green = 8'h97;    Blue = 8'h5d;
end 13'h1698:    begin Red = 8'h71;    Green = 8'h52;    Blue = 8'h26;
end 13'h1699:    begin Red = 8'hb3;    Green = 8'h81;    Blue = 8'h4c;
end 13'h169a:    begin Red = 8'hb0;    Green = 8'h82;    Blue = 8'h50;
end 13'h169b:    begin Red = 8'haf;    Green = 8'h85;    Blue = 8'h49;
end 13'h169c:    begin Red = 8'haa;    Green = 8'h83;    Blue = 8'h4c;
end 13'h169d:    begin Red = 8'h70;    Green = 8'h5a;    Blue = 8'h2b;
end 13'h169e:    begin Red = 8'h94;    Green = 8'h72;    Blue = 8'h44;
end 13'h169f:    begin Red = 8'h8a;    Green = 8'h64;    Blue = 8'h40;
end 13'h16a0:    begin Red = 8'hca;    Green = 8'hc3;    Blue = 8'h9b;
end 13'h16a1:    begin Red = 8'h00;    Green = 8'h53;    Blue = 8'h10;
end 13'h16a2:    begin Red = 8'h35;    Green = 8'h29;    Blue = 8'h2d;
end 13'h16a3:    begin Red = 8'h31;    Green = 8'h28;    Blue = 8'h29;
end 13'h16a4:    begin Red = 8'h2f;    Green = 8'h2a;    Blue = 8'h27;
end 13'h16a5:    begin Red = 8'h3a;    Green = 8'h30;    Blue = 8'h2e;
end 13'h16a6:    begin Red = 8'h3b;    Green = 8'h2f;    Blue = 8'h33;
end 13'h16a7:    begin Red = 8'h00;    Green = 8'hfc;    Blue = 8'h17;
end 13'h16a8:    begin Red = 8'heb;    Green = 8'hea;    Blue = 8'hda;
end 13'h16a9:    begin Red = 8'hfa;    Green = 8'hf1;    Blue = 8'he4;
end 13'h16aa:    begin Red = 8'ha3;    Green = 8'h7d;    Blue = 8'h61;
end 13'h16ab:    begin Red = 8'h97;    Green = 8'h88;    Blue = 8'h5b;
end 13'h16ac:    begin Red = 8'h9a;    Green = 8'h90;    Blue = 8'h5a;
end 13'h16ad:    begin Red = 8'h7a;    Green = 8'h75;    Blue = 8'h53;
end 13'h16ae:    begin Red = 8'h63;    Green = 8'h66;    Blue = 8'h3f;
end 13'h16af:    begin Red = 8'hb9;    Green = 8'hb8;    Blue = 8'h94;
end 13'h16b0:    begin Red = 8'h87;    Green = 8'h72;    Blue = 8'h56;
end 13'h16b1:    begin Red = 8'h88;    Green = 8'h74;    Blue = 8'h58;
end 13'h16b2:    begin Red = 8'h6e;    Green = 8'h67;    Blue = 8'h45;
end 13'h16b3:    begin Red = 8'h6f;    Green = 8'h53;    Blue = 8'h2c;
end 13'h16b4:    begin Red = 8'h82;    Green = 8'h61;    Blue = 8'h36;
end 13'h16b5:    begin Red = 8'hba;    Green = 8'h92;    Blue = 8'h55;
end 13'h16b6:    begin Red = 8'ha3;    Green = 8'h7b;    Blue = 8'h47;
end 13'h16b7:    begin Red = 8'h9d;    Green = 8'h7c;    Blue = 8'h47;
end 13'h16b8:    begin Red = 8'h9f;    Green = 8'h79;    Blue = 8'h48;
end 13'h16b9:    begin Red = 8'hc0;    Green = 8'hcd;    Blue = 8'hb0;
end 13'h16ba:    begin Red = 8'h99;    Green = 8'h73;    Blue = 8'h42;
end 13'h16bb:    begin Red = 8'h8a;    Green = 8'h77;    Blue = 8'h57;
end 13'h16bc:    begin Red = 8'h9c;    Green = 8'h8a;    Blue = 8'h5a;
end 13'h16bd:    begin Red = 8'h00;    Green = 8'h05;    Blue = 8'h05;
end 13'h16be:    begin Red = 8'h33;    Green = 8'h28;    Blue = 8'h26;
end 13'h16bf:    begin Red = 8'h31;    Green = 8'h26;    Blue = 8'h24;
end 13'h16c0:    begin Red = 8'h40;    Green = 8'h31;    Blue = 8'h2c;
end 13'h16c1:    begin Red = 8'h01;    Green = 8'h5f;    Blue = 8'h13;
end 13'h16c2:    begin Red = 8'h2c;    Green = 8'h22;    Blue = 8'h19;
end 13'h16c3:    begin Red = 8'h34;    Green = 8'h22;    Blue = 8'h18;
end 13'h16c4:    begin Red = 8'h2f;    Green = 8'h21;    Blue = 8'h18;
end 13'h16c5:    begin Red = 8'h32;    Green = 8'h1f;    Blue = 8'h18;
end 13'h16c6:    begin Red = 8'h30;    Green = 8'h1c;    Blue = 8'h15;
end 13'h16c7:    begin Red = 8'h2b;    Green = 8'h22;    Blue = 8'h11;
end 13'h16c8:    begin Red = 8'h38;    Green = 8'h1f;    Blue = 8'h1a;
end 13'h16c9:    begin Red = 8'h03;    Green = 8'h52;    Blue = 8'h19;
end 13'h16ca:    begin Red = 8'h37;    Green = 8'h21;    Blue = 8'h13;
end 13'h16cb:    begin Red = 8'h2e;    Green = 8'h20;    Blue = 8'h15;
end 13'h16cc:    begin Red = 8'h35;    Green = 8'h1d;    Blue = 8'h19;
end 13'h16cd:    begin Red = 8'h00;    Green = 8'h01;    Blue = 8'h32;
end 13'h16ce:    begin Red = 8'hd4;    Green = 8'hb6;    Blue = 8'h90;
end 13'h16cf:    begin Red = 8'h4e;    Green = 8'h4f;    Blue = 8'h53;
end 13'h16d0:    begin Red = 8'h4f;    Green = 8'h50;    Blue = 8'h4a;
end 13'h16d1:    begin Red = 8'h4d;    Green = 8'h4e;    Blue = 8'h48;
end 13'h16d2:    begin Red = 8'hf6;    Green = 8'hf3;    Blue = 8'hc0;
end 13'h16d3:    begin Red = 8'hf9;    Green = 8'hd3;    Blue = 8'ha2;
end 13'h16d4:    begin Red = 8'he2;    Green = 8'hc8;    Blue = 8'h9e;
end 13'h16d5:    begin Red = 8'hde;    Green = 8'hcd;    Blue = 8'hb6;
end 13'h16d6:    begin Red = 8'hf2;    Green = 8'he6;    Blue = 8'hd4;
end 13'h16d7:    begin Red = 8'h49;    Green = 8'h41;    Blue = 8'h48;
end 13'h16d8:    begin Red = 8'he7;    Green = 8'hd6;    Blue = 8'hc3;
end 13'h16d9:    begin Red = 8'hb1;    Green = 8'hae;    Blue = 8'h74;
end 13'h16da:    begin Red = 8'h91;    Green = 8'h8a;    Blue = 8'h56;
end 13'h16db:    begin Red = 8'h97;    Green = 8'h8d;    Blue = 8'h5d;
end 13'h16dc:    begin Red = 8'h70;    Green = 8'h71;    Blue = 8'h72;
end 13'h16dd:    begin Red = 8'h73;    Green = 8'h70;    Blue = 8'h6d;
end 13'h16de:    begin Red = 8'h74;    Green = 8'h78;    Blue = 8'h72;
end 13'h16df:    begin Red = 8'h6f;    Green = 8'h76;    Blue = 8'h65;
end 13'h16e0:    begin Red = 8'h7d;    Green = 8'h70;    Blue = 8'h72;
end 13'h16e1:    begin Red = 8'he9;    Green = 8'he2;    Blue = 8'hc7;
end 13'h16e2:    begin Red = 8'hc8;    Green = 8'hba;    Blue = 8'ha7;
end 13'h16e3:    begin Red = 8'hbe;    Green = 8'hc2;    Blue = 8'h97;
end 13'h16e4:    begin Red = 8'h7b;    Green = 8'h68;    Blue = 8'h4a;
end 13'h16e5:    begin Red = 8'h04;    Green = 8'h21;    Blue = 8'hb0;
end 13'h16e6:    begin Red = 8'h05;    Green = 8'he3;    Blue = 8'h94;
end 13'h16e7:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'h39;
end 13'h16e8:    begin Red = 8'h08;    Green = 8'h65;    Blue = 8'h4d;
end 13'h16e9:    begin Red = 8'h08;    Green = 8'h04;    Blue = 8'hdb;
end 13'h16ea:    begin Red = 8'h7e;    Green = 8'h4e;    Blue = 8'h10;
end 13'h16eb:    begin Red = 8'h07;    Green = 8'he4;    Blue = 8'hec;
end 13'h16ec:    begin Red = 8'h07;    Green = 8'hf4;    Blue = 8'hfd;
end 13'h16ed:    begin Red = 8'h07;    Green = 8'he4;    Blue = 8'hfb;
end 13'h16ee:    begin Red = 8'h07;    Green = 8'hb5;    Blue = 8'h0c;
end 13'h16ef:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h35;
end 13'h16f0:    begin Red = 8'h05;    Green = 8'h83;    Blue = 8'h39;
end 13'h16f1:    begin Red = 8'h05;    Green = 8'h33;    Blue = 8'h06;
end 13'h16f2:    begin Red = 8'h07;    Green = 8'hb4;    Blue = 8'h7d;
end 13'h16f3:    begin Red = 8'h07;    Green = 8'h34;    Blue = 8'h6f;
end 13'h16f4:    begin Red = 8'h07;    Green = 8'h14;    Blue = 8'h4b;
end 13'h16f5:    begin Red = 8'h06;    Green = 8'hf4;    Blue = 8'h5b;
end 13'h16f6:    begin Red = 8'h07;    Green = 8'h04;    Blue = 8'h6c;
end 13'h16f7:    begin Red = 8'he7;    Green = 8'hf3;    Blue = 8'hd4;
end 13'h16f8:    begin Red = 8'h67;    Green = 8'h47;    Blue = 8'h16;
end 13'h16f9:    begin Red = 8'h6a;    Green = 8'h49;    Blue = 8'h13;
end 13'h16fa:    begin Red = 8'h06;    Green = 8'h84;    Blue = 8'h4a;
end 13'h16fb:    begin Red = 8'h05;    Green = 8'hf3;    Blue = 8'hdd;
end 13'h16fc:    begin Red = 8'ha0;    Green = 8'ha6;    Blue = 8'h8d;
end 13'h16fd:    begin Red = 8'h8f;    Green = 8'h74;    Blue = 8'h59;
end 13'h16fe:    begin Red = 8'h29;    Green = 8'h1d;    Blue = 8'h1f;
end 13'h16ff:    begin Red = 8'h34;    Green = 8'h25;    Blue = 8'h22;
end 13'h1700:    begin Red = 8'h00;    Green = 8'h0a;    Blue = 8'h46;
end 13'h1701:    begin Red = 8'h2b;    Green = 8'h1e;    Blue = 8'h16;
end 13'h1702:    begin Red = 8'h02;    Green = 8'h61;    Blue = 8'he9;
end 13'h1703:    begin Red = 8'h1f;    Green = 8'h1a;    Blue = 8'h16;
end 13'h1704:    begin Red = 8'h02;    Green = 8'h91;    Blue = 8'hec;
end 13'h1705:    begin Red = 8'h39;    Green = 8'h25;    Blue = 8'h1e;
end 13'h1706:    begin Red = 8'h38;    Green = 8'h27;    Blue = 8'h20;
end 13'h1707:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'hbb;
end 13'h1708:    begin Red = 8'h02;    Green = 8'h31;    Blue = 8'he1;
end 13'h1709:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'hdd;
end 13'h170a:    begin Red = 8'h02;    Green = 8'h41;    Blue = 8'h93;
end 13'h170b:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'hff;
end 13'h170c:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'hfd;
end 13'h170d:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'hca;
end 13'h170e:    begin Red = 8'h02;    Green = 8'h62;    Blue = 8'h06;
end 13'h170f:    begin Red = 8'h36;    Green = 8'h22;    Blue = 8'h1b;
end 13'h1710:    begin Red = 8'h2b;    Green = 8'h1d;    Blue = 8'h10;
end 13'h1711:    begin Red = 8'h00;    Green = 8'h08;    Blue = 8'h02;
end 13'h1712:    begin Red = 8'hee;    Green = 8'hdc;    Blue = 8'hac;
end 13'h1713:    begin Red = 8'hef;    Green = 8'hc5;    Blue = 8'h95;
end 13'h1714:    begin Red = 8'hfb;    Green = 8'hd7;    Blue = 8'h99;
end 13'h1715:    begin Red = 8'h47;    Green = 8'h4e;    Blue = 8'h56;
end 13'h1716:    begin Red = 8'h2b;    Green = 8'h35;    Blue = 8'h50;
end 13'h1717:    begin Red = 8'h33;    Green = 8'h3a;    Blue = 8'h56;
end 13'h1718:    begin Red = 8'h9b;    Green = 8'h9b;    Blue = 8'h72;
end 13'h1719:    begin Red = 8'hd2;    Green = 8'hde;    Blue = 8'hca;
end 13'h171a:    begin Red = 8'hd6;    Green = 8'he0;    Blue = 8'hcd;
end 13'h171b:    begin Red = 8'hf9;    Green = 8'hff;    Blue = 8'hed;
end 13'h171c:    begin Red = 8'hfa;    Green = 8'hf2;    Blue = 8'hea;
end 13'h171d:    begin Red = 8'h45;    Green = 8'h42;    Blue = 8'h4a;
end 13'h171e:    begin Red = 8'h46;    Green = 8'h3d;    Blue = 8'h42;
end 13'h171f:    begin Red = 8'hb2;    Green = 8'hb2;    Blue = 8'h62;
end 13'h1720:    begin Red = 8'h97;    Green = 8'h8a;    Blue = 8'h63;
end 13'h1721:    begin Red = 8'h5d;    Green = 8'h5c;    Blue = 8'h75;
end 13'h1722:    begin Red = 8'h64;    Green = 8'h61;    Blue = 8'h77;
end 13'h1723:    begin Red = 8'h65;    Green = 8'h5e;    Blue = 8'h74;
end 13'h1724:    begin Red = 8'h77;    Green = 8'h72;    Blue = 8'h75;
end 13'h1725:    begin Red = 8'hd7;    Green = 8'hd2;    Blue = 8'hbb;
end 13'h1726:    begin Red = 8'hdd;    Green = 8'he2;    Blue = 8'hc5;
end 13'h1727:    begin Red = 8'h6f;    Green = 8'h5d;    Blue = 8'h34;
end 13'h1728:    begin Red = 8'h68;    Green = 8'h53;    Blue = 8'h36;
end 13'h1729:    begin Red = 8'h04;    Green = 8'h01;    Blue = 8'he3;
end 13'h172a:    begin Red = 8'h05;    Green = 8'hd3;    Blue = 8'h54;
end 13'h172b:    begin Red = 8'h08;    Green = 8'hd5;    Blue = 8'h7d;
end 13'h172c:    begin Red = 8'h08;    Green = 8'h75;    Blue = 8'h2c;
end 13'h172d:    begin Red = 8'h84;    Green = 8'h51;    Blue = 8'h10;
end 13'h172e:    begin Red = 8'h08;    Green = 8'h45;    Blue = 8'h1f;
end 13'h172f:    begin Red = 8'h08;    Green = 8'h35;    Blue = 8'h3b;
end 13'h1730:    begin Red = 8'h08;    Green = 8'h15;    Blue = 8'h0d;
end 13'h1731:    begin Red = 8'he8;    Green = 8'hb5;    Blue = 8'h7c;
end 13'h1732:    begin Red = 8'h05;    Green = 8'h63;    Blue = 8'h6d;
end 13'h1733:    begin Red = 8'h05;    Green = 8'h93;    Blue = 8'h47;
end 13'h1734:    begin Red = 8'h05;    Green = 8'h63;    Blue = 8'h46;
end 13'h1735:    begin Red = 8'h07;    Green = 8'hd4;    Blue = 8'hdd;
end 13'h1736:    begin Red = 8'h07;    Green = 8'h14;    Blue = 8'h8a;
end 13'h1737:    begin Red = 8'h07;    Green = 8'h14;    Blue = 8'h9b;
end 13'h1738:    begin Red = 8'h07;    Green = 8'h04;    Blue = 8'h8b;
end 13'h1739:    begin Red = 8'he0;    Green = 8'hed;    Blue = 8'hd0;
end 13'h173a:    begin Red = 8'h6b;    Green = 8'h46;    Blue = 8'h12;
end 13'h173b:    begin Red = 8'h06;    Green = 8'hc4;    Blue = 8'h5c;
end 13'h173c:    begin Red = 8'h06;    Green = 8'ha4;    Blue = 8'h25;
end 13'h173d:    begin Red = 8'h06;    Green = 8'h23;    Blue = 8'hd8;
end 13'h173e:    begin Red = 8'hdc;    Green = 8'hd4;    Blue = 8'had;
end 13'h173f:    begin Red = 8'h8b;    Green = 8'h68;    Blue = 8'h17;
end 13'h1740:    begin Red = 8'h92;    Green = 8'h67;    Blue = 8'h19;
end 13'h1741:    begin Red = 8'h85;    Green = 8'h6b;    Blue = 8'h17;
end 13'h1742:    begin Red = 8'h8a;    Green = 8'h6b;    Blue = 8'h11;
end 13'h1743:    begin Red = 8'h07;    Green = 8'hf6;    Blue = 8'hc5;
end 13'h1744:    begin Red = 8'h08;    Green = 8'h46;    Blue = 8'h36;
end 13'h1745:    begin Red = 8'h3f;    Green = 8'h35;    Blue = 8'h29;
end 13'h1746:    begin Red = 8'hff;    Green = 8'hfa;    Blue = 8'hc3;
end 13'h1747:    begin Red = 8'h4c;    Green = 8'h34;    Blue = 8'h34;
end 13'h1748:    begin Red = 8'h41;    Green = 8'h2c;    Blue = 8'h29;
end 13'h1749:    begin Red = 8'h42;    Green = 8'h28;    Blue = 8'h2b;
end 13'h174a:    begin Red = 8'h21;    Green = 8'h16;    Blue = 8'h10;
end 13'h174b:    begin Red = 8'h00;    Green = 8'h14;    Blue = 8'he2;
end 13'h174c:    begin Red = 8'h4b;    Green = 8'h30;    Blue = 8'h35;
end 13'h174d:    begin Red = 8'h48;    Green = 8'h2f;    Blue = 8'h32;
end 13'h174e:    begin Red = 8'h71;    Green = 8'h3d;    Blue = 8'h64;
end 13'h174f:    begin Red = 8'h66;    Green = 8'h39;    Blue = 8'h56;
end 13'h1750:    begin Red = 8'h5d;    Green = 8'h37;    Blue = 8'h5c;
end 13'h1751:    begin Red = 8'h38;    Green = 8'h26;    Blue = 8'h24;
end 13'h1752:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h4e;
end 13'h1753:    begin Red = 8'h00;    Green = 8'h14;    Blue = 8'hd7;
end 13'h1754:    begin Red = 8'h4c;    Green = 8'h31;    Blue = 8'h38;
end 13'h1755:    begin Red = 8'h46;    Green = 8'h2d;    Blue = 8'h30;
end 13'h1756:    begin Red = 8'h44;    Green = 8'h2b;    Blue = 8'h31;
end 13'h1757:    begin Red = 8'h41;    Green = 8'h2b;    Blue = 8'h2d;
end 13'h1758:    begin Red = 8'h3d;    Green = 8'h29;    Blue = 8'h2b;
end 13'h1759:    begin Red = 8'h00;    Green = 8'h13;    Blue = 8'h0d;
end 13'h175a:    begin Red = 8'h2d;    Green = 8'h2e;    Blue = 8'h33;
end 13'h175b:    begin Red = 8'h2d;    Green = 8'h26;    Blue = 8'h20;
end 13'h175c:    begin Red = 8'h00;    Green = 8'h95;    Blue = 8'h1c;
end 13'h175d:    begin Red = 8'hd3;    Green = 8'ha7;    Blue = 8'h24;
end 13'h175e:    begin Red = 8'h51;    Green = 8'h53;    Blue = 8'h48;
end 13'h175f:    begin Red = 8'hc7;    Green = 8'h67;    Blue = 8'h61;
end 13'h1760:    begin Red = 8'he5;    Green = 8'hd3;    Blue = 8'hbb;
end 13'h1761:    begin Red = 8'h57;    Green = 8'h50;    Blue = 8'h52;
end 13'h1762:    begin Red = 8'h5a;    Green = 8'h51;    Blue = 8'h59;
end 13'h1763:    begin Red = 8'h46;    Green = 8'h3e;    Blue = 8'h46;
end 13'h1764:    begin Red = 8'hae;    Green = 8'hb3;    Blue = 8'h66;
end 13'h1765:    begin Red = 8'h8d;    Green = 8'h80;    Blue = 8'h5a;
end 13'h1766:    begin Red = 8'h9a;    Green = 8'h8e;    Blue = 8'h57;
end 13'h1767:    begin Red = 8'h72;    Green = 8'h73;    Blue = 8'h6e;
end 13'h1768:    begin Red = 8'h7a;    Green = 8'h7b;    Blue = 8'h76;
end 13'h1769:    begin Red = 8'hdb;    Green = 8'hb9;    Blue = 8'h51;
end 13'h176a:    begin Red = 8'hde;    Green = 8'hb8;    Blue = 8'h4f;
end 13'h176b:    begin Red = 8'h38;    Green = 8'h39;    Blue = 8'h49;
end 13'h176c:    begin Red = 8'h75;    Green = 8'h75;    Blue = 8'h6e;
end 13'h176d:    begin Red = 8'h75;    Green = 8'h75;    Blue = 8'h77;
end 13'h176e:    begin Red = 8'h02;    Green = 8'hf1;    Blue = 8'h40;
end 13'h176f:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'he1;
end 13'h1770:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'hb2;
end 13'h1771:    begin Red = 8'h06;    Green = 8'hb4;    Blue = 8'h38;
end 13'h1772:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'hf4;
end 13'h1773:    begin Red = 8'h06;    Green = 8'hd4;    Blue = 8'h14;
end 13'h1774:    begin Red = 8'h06;    Green = 8'hc4;    Blue = 8'h03;
end 13'h1775:    begin Red = 8'h06;    Green = 8'h93;    Blue = 8'hf5;
end 13'h1776:    begin Red = 8'h06;    Green = 8'ha4;    Blue = 8'h06;
end 13'h1777:    begin Red = 8'h06;    Green = 8'h84;    Blue = 8'h16;
end 13'h1778:    begin Red = 8'h06;    Green = 8'h63;    Blue = 8'hf4;
end 13'h1779:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'hdb;
end 13'h177a:    begin Red = 8'h04;    Green = 8'h42;    Blue = 8'h81;
end 13'h177b:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h60;
end 13'h177c:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h91;
end 13'h177d:    begin Red = 8'h06;    Green = 8'h03;    Blue = 8'hf9;
end 13'h177e:    begin Red = 8'h05;    Green = 8'hd3;    Blue = 8'hd4;
end 13'h177f:    begin Red = 8'h05;    Green = 8'hf3;    Blue = 8'hc4;
end 13'h1780:    begin Red = 8'h05;    Green = 8'h93;    Blue = 8'h83;
end 13'h1781:    begin Red = 8'heb;    Green = 8'hf0;    Blue = 8'hd3;
end 13'h1782:    begin Red = 8'h05;    Green = 8'h73;    Blue = 8'h58;
end 13'h1783:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h25;
end 13'h1784:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h56;
end 13'h1785:    begin Red = 8'h05;    Green = 8'h23;    Blue = 8'h23;
end 13'h1786:    begin Red = 8'h05;    Green = 8'h33;    Blue = 8'h14;
end 13'h1787:    begin Red = 8'h04;    Green = 8'he3;    Blue = 8'h87;
end 13'h1788:    begin Red = 8'h33;    Green = 8'h40;    Blue = 8'h75;
end 13'h1789:    begin Red = 8'h30;    Green = 8'h46;    Blue = 8'h6f;
end 13'h178a:    begin Red = 8'h2c;    Green = 8'h48;    Blue = 8'h6f;
end 13'h178b:    begin Red = 8'h81;    Green = 8'h6b;    Blue = 8'h15;
end 13'h178c:    begin Red = 8'hc0;    Green = 8'hab;    Blue = 8'h76;
end 13'h178d:    begin Red = 8'hc4;    Green = 8'haa;    Blue = 8'h79;
end 13'h178e:    begin Red = 8'hc4;    Green = 8'hab;    Blue = 8'h73;
end 13'h178f:    begin Red = 8'hc0;    Green = 8'ha8;    Blue = 8'h78;
end 13'h1790:    begin Red = 8'h50;    Green = 8'h3a;    Blue = 8'h3c;
end 13'h1791:    begin Red = 8'h4e;    Green = 8'h32;    Blue = 8'h40;
end 13'h1792:    begin Red = 8'h4d;    Green = 8'h36;    Blue = 8'h40;
end 13'h1793:    begin Red = 8'h01;    Green = 8'hf1;    Blue = 8'h4e;
end 13'h1794:    begin Red = 8'h59;    Green = 8'h3e;    Blue = 8'h47;
end 13'h1795:    begin Red = 8'h55;    Green = 8'h3c;    Blue = 8'h42;
end 13'h1796:    begin Red = 8'h58;    Green = 8'h3a;    Blue = 8'h46;
end 13'h1797:    begin Red = 8'h47;    Green = 8'h2d;    Blue = 8'h36;
end 13'h1798:    begin Red = 8'h46;    Green = 8'h36;    Blue = 8'h36;
end 13'h1799:    begin Red = 8'h4a;    Green = 8'h35;    Blue = 8'h3a;
end 13'h179a:    begin Red = 8'h43;    Green = 8'h34;    Blue = 8'h3b;
end 13'h179b:    begin Red = 8'h4b;    Green = 8'h38;    Blue = 8'h3c;
end 13'h179c:    begin Red = 8'h4e;    Green = 8'h33;    Blue = 8'h3c;
end 13'h179d:    begin Red = 8'h3f;    Green = 8'h2c;    Blue = 8'h30;
end 13'h179e:    begin Red = 8'h41;    Green = 8'h2b;    Blue = 8'h38;
end 13'h179f:    begin Red = 8'h44;    Green = 8'h31;    Blue = 8'h37;
end 13'h17a0:    begin Red = 8'h01;    Green = 8'h6d;    Blue = 8'h10;
end 13'h17a1:    begin Red = 8'h5b;    Green = 8'h3f;    Blue = 8'h4e;
end 13'h17a2:    begin Red = 8'h56;    Green = 8'h3b;    Blue = 8'h4a;
end 13'h17a3:    begin Red = 8'h53;    Green = 8'h38;    Blue = 8'h49;
end 13'h17a4:    begin Red = 8'h50;    Green = 8'h35;    Blue = 8'h46;
end 13'h17a5:    begin Red = 8'h4b;    Green = 8'h33;    Blue = 8'h41;
end 13'h17a6:    begin Red = 8'h02;    Green = 8'h2b;    Blue = 8'h25;
end 13'h17a7:    begin Red = 8'hf3;    Green = 8'hef;    Blue = 8'hde;
end 13'h17a8:    begin Red = 8'hca;    Green = 8'hbb;    Blue = 8'h71;
end 13'h17a9:    begin Red = 8'hf5;    Green = 8'hef;    Blue = 8'hea;
end 13'h17aa:    begin Red = 8'hc3;    Green = 8'haf;    Blue = 8'h6b;
end 13'h17ab:    begin Red = 8'h34;    Green = 8'h58;    Blue = 8'h84;
end 13'h17ac:    begin Red = 8'h3f;    Green = 8'h61;    Blue = 8'h7d;
end 13'h17ad:    begin Red = 8'h39;    Green = 8'h61;    Blue = 8'h7e;
end 13'h17ae:    begin Red = 8'h3f;    Green = 8'h68;    Blue = 8'h85;
end 13'h17af:    begin Red = 8'h75;    Green = 8'hce;    Blue = 8'hff;
end 13'h17b0:    begin Red = 8'h72;    Green = 8'hcc;    Blue = 8'hff;
end 13'h17b1:    begin Red = 8'hdf;    Green = 8'hff;    Blue = 8'hff;
end 13'h17b2:    begin Red = 8'hde;    Green = 8'hfe;    Blue = 8'hf7;
end 13'h17b3:    begin Red = 8'hcc;    Green = 8'h77;    Blue = 8'h7c;
end 13'h17b4:    begin Red = 8'hbb;    Green = 8'hc1;    Blue = 8'h98;
end 13'h17b5:    begin Red = 8'h04;    Green = 8'he2;    Blue = 8'hc6;
end 13'h17b6:    begin Red = 8'hb1;    Green = 8'hae;    Blue = 8'h7b;
end 13'h17b7:    begin Red = 8'ha6;    Green = 8'ha5;    Blue = 8'h75;
end 13'h17b8:    begin Red = 8'ha1;    Green = 8'ha4;    Blue = 8'h6f;
end 13'h17b9:    begin Red = 8'h9b;    Green = 8'ha2;    Blue = 8'h6c;
end 13'h17ba:    begin Red = 8'h96;    Green = 8'h95;    Blue = 8'h65;
end 13'h17bb:    begin Red = 8'h9c;    Green = 8'h9b;    Blue = 8'h6b;
end 13'h17bc:    begin Red = 8'h88;    Green = 8'h91;    Blue = 8'h62;
end 13'h17bd:    begin Red = 8'h75;    Green = 8'h83;    Blue = 8'h4e;
end 13'h17be:    begin Red = 8'h06;    Green = 8'h83;    Blue = 8'h61;
end 13'h17bf:    begin Red = 8'hee;    Green = 8'hbe;    Blue = 8'h80;
end 13'h17c0:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'h77;
end 13'h17c1:    begin Red = 8'h99;    Green = 8'h9a;    Blue = 8'h6e;
end 13'h17c2:    begin Red = 8'h93;    Green = 8'h90;    Blue = 8'h67;
end 13'h17c3:    begin Red = 8'h8e;    Green = 8'h8f;    Blue = 8'h63;
end 13'h17c4:    begin Red = 8'h86;    Green = 8'h8c;    Blue = 8'h5c;
end 13'h17c5:    begin Red = 8'hc3;    Green = 8'hcc;    Blue = 8'hac;
end 13'h17c6:    begin Red = 8'h4d;    Green = 8'h5f;    Blue = 8'h37;
end 13'h17c7:    begin Red = 8'h47;    Green = 8'h59;    Blue = 8'h2f;
end 13'h17c8:    begin Red = 8'h05;    Green = 8'h23;    Blue = 8'hac;
end 13'h17c9:    begin Red = 8'h15;    Green = 8'h2b;    Blue = 8'h39;
end 13'h17ca:    begin Red = 8'h17;    Green = 8'h29;    Blue = 8'h3f;
end 13'h17cb:    begin Red = 8'h20;    Green = 8'h2c;    Blue = 8'h44;
end 13'h17cc:    begin Red = 8'h2d;    Green = 8'h2d;    Blue = 8'h47;
end 13'h17cd:    begin Red = 8'h2c;    Green = 8'h31;    Blue = 8'h44;
end 13'h17ce:    begin Red = 8'h3f;    Green = 8'h4f;    Blue = 8'h5e;
end 13'h17cf:    begin Red = 8'h3f;    Green = 8'h45;    Blue = 8'h53;
end 13'h17d0:    begin Red = 8'h3d;    Green = 8'h40;    Blue = 8'h51;
end 13'h17d1:    begin Red = 8'h39;    Green = 8'h45;    Blue = 8'h5b;
end 13'h17d2:    begin Red = 8'h3a;    Green = 8'h49;    Blue = 8'h60;
end 13'h17d3:    begin Red = 8'h37;    Green = 8'h46;    Blue = 8'h49;
end 13'h17d4:    begin Red = 8'h37;    Green = 8'h44;    Blue = 8'h55;
end 13'h17d5:    begin Red = 8'h3b;    Green = 8'h41;    Blue = 8'h4d;
end 13'h17d6:    begin Red = 8'h88;    Green = 8'h6d;    Blue = 8'h16;
end 13'h17d7:    begin Red = 8'h08;    Green = 8'h26;    Blue = 8'h36;
end 13'h17d8:    begin Red = 8'had;    Green = 8'h94;    Blue = 8'h80;
end 13'h17d9:    begin Red = 8'hca;    Green = 8'hb3;    Blue = 8'h7f;
end 13'h17da:    begin Red = 8'hcf;    Green = 8'hb6;    Blue = 8'h7e;
end 13'h17db:    begin Red = 8'hd1;    Green = 8'hb8;    Blue = 8'h80;
end 13'h17dc:    begin Red = 8'hba;    Green = 8'ha0;    Blue = 8'h6f;
end 13'h17dd:    begin Red = 8'h48;    Green = 8'h32;    Blue = 8'h34;
end 13'h17de:    begin Red = 8'h4f;    Green = 8'h38;    Blue = 8'h42;
end 13'h17df:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h7d;
end 13'h17e0:    begin Red = 8'h5a;    Green = 8'h40;    Blue = 8'h49;
end 13'h17e1:    begin Red = 8'h58;    Green = 8'h38;    Blue = 8'h43;
end 13'h17e2:    begin Red = 8'h4d;    Green = 8'h3e;    Blue = 8'h43;
end 13'h17e3:    begin Red = 8'h47;    Green = 8'h2c;    Blue = 8'h3b;
end 13'h17e4:    begin Red = 8'h4d;    Green = 8'h2e;    Blue = 8'h3d;
end 13'h17e5:    begin Red = 8'h52;    Green = 8'h33;    Blue = 8'h45;
end 13'h17e6:    begin Red = 8'h43;    Green = 8'h2c;    Blue = 8'h40;
end 13'h17e7:    begin Red = 8'h43;    Green = 8'h31;    Blue = 8'h3f;
end 13'h17e8:    begin Red = 8'h45;    Green = 8'h35;    Blue = 8'h40;
end 13'h17e9:    begin Red = 8'h45;    Green = 8'h30;    Blue = 8'h43;
end 13'h17ea:    begin Red = 8'h02;    Green = 8'h01;    Blue = 8'h76;
end 13'h17eb:    begin Red = 8'h00;    Green = 8'h11;    Blue = 8'hd4;
end 13'h17ec:    begin Red = 8'h4f;    Green = 8'h35;    Blue = 8'h3e;
end 13'h17ed:    begin Red = 8'h51;    Green = 8'h39;    Blue = 8'h46;
end 13'h17ee:    begin Red = 8'h1c;    Green = 8'h10;    Blue = 8'h1c;
end 13'h17ef:    begin Red = 8'hc5;    Green = 8'h67;    Blue = 8'h65;
end 13'h17f0:    begin Red = 8'hc9;    Green = 8'h68;    Blue = 8'h64;
end 13'h17f1:    begin Red = 8'hc6;    Green = 8'h68;    Blue = 8'h5e;
end 13'h17f2:    begin Red = 8'hca;    Green = 8'hc0;    Blue = 8'h6f;
end 13'h17f3:    begin Red = 8'hbd;    Green = 8'h9b;    Blue = 8'h57;
end 13'h17f4:    begin Red = 8'hc7;    Green = 8'ha8;    Blue = 8'h69;
end 13'h17f5:    begin Red = 8'h43;    Green = 8'h6b;    Blue = 8'h7d;
end 13'h17f6:    begin Red = 8'h56;    Green = 8'h7d;    Blue = 8'h95;
end 13'h17f7:    begin Red = 8'h5d;    Green = 8'h7d;    Blue = 8'h98;
end 13'h17f8:    begin Red = 8'h4c;    Green = 8'h80;    Blue = 8'h94;
end 13'h17f9:    begin Red = 8'h74;    Green = 8'hd9;    Blue = 8'hf6;
end 13'h17fa:    begin Red = 8'h75;    Green = 8'hb6;    Blue = 8'he2;
end 13'h17fb:    begin Red = 8'h73;    Green = 8'hbe;    Blue = 8'hf1;
end 13'h17fc:    begin Red = 8'hd9;    Green = 8'hf3;    Blue = 8'hfd;
end 13'h17fd:    begin Red = 8'he2;    Green = 8'hfd;    Blue = 8'hf8;
end 13'h17fe:    begin Red = 8'hde;    Green = 8'h74;    Blue = 8'h66;
end 13'h17ff:    begin Red = 8'hed;    Green = 8'hf1;    Blue = 8'hc7;
end 13'h1800:    begin Red = 8'h9d;    Green = 8'h8b;    Blue = 8'h53;
end 13'h1801:    begin Red = 8'h95;    Green = 8'h86;    Blue = 8'h58;
end 13'h1802:    begin Red = 8'h9b;    Green = 8'h86;    Blue = 8'h5a;
end 13'h1803:    begin Red = 8'h9c;    Green = 8'h91;    Blue = 8'h55;
end 13'h1804:    begin Red = 8'h34;    Green = 8'h34;    Blue = 8'h48;
end 13'h1805:    begin Red = 8'hc8;    Green = 8'hbb;    Blue = 8'haf;
end 13'h1806:    begin Red = 8'he6;    Green = 8'hbd;    Blue = 8'h7b;
end 13'h1807:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'he2;
end 13'h1808:    begin Red = 8'h6f;    Green = 8'h69;    Blue = 8'h47;
end 13'h1809:    begin Red = 8'ha4;    Green = 8'h9e;    Blue = 8'h6a;
end 13'h180a:    begin Red = 8'h9c;    Green = 8'h94;    Blue = 8'h65;
end 13'h180b:    begin Red = 8'h97;    Green = 8'h92;    Blue = 8'h5b;
end 13'h180c:    begin Red = 8'h98;    Green = 8'h92;    Blue = 8'h60;
end 13'h180d:    begin Red = 8'h94;    Green = 8'h91;    Blue = 8'h5e;
end 13'h180e:    begin Red = 8'h85;    Green = 8'h83;    Blue = 8'h53;
end 13'h180f:    begin Red = 8'h61;    Green = 8'h68;    Blue = 8'h3c;
end 13'h1810:    begin Red = 8'h5b;    Green = 8'h67;    Blue = 8'h39;
end 13'h1811:    begin Red = 8'h06;    Green = 8'h13;    Blue = 8'hd3;
end 13'h1812:    begin Red = 8'hda;    Green = 8'hb3;    Blue = 8'h72;
end 13'h1813:    begin Red = 8'hb7;    Green = 8'hc1;    Blue = 8'h9f;
end 13'h1814:    begin Red = 8'h5c;    Green = 8'h61;    Blue = 8'h38;
end 13'h1815:    begin Red = 8'h52;    Green = 8'h57;    Blue = 8'h2e;
end 13'h1816:    begin Red = 8'h4b;    Green = 8'h52;    Blue = 8'h28;
end 13'h1817:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h88;
end 13'h1818:    begin Red = 8'hac;    Green = 8'h8a;    Blue = 8'h5a;
end 13'h1819:    begin Red = 8'h86;    Green = 8'h65;    Blue = 8'h3a;
end 13'h181a:    begin Red = 8'h6b;    Green = 8'hc9;    Blue = 8'hd3;
end 13'h181b:    begin Red = 8'h81;    Green = 8'hd1;    Blue = 8'hce;
end 13'h181c:    begin Red = 8'h3a;    Green = 8'h51;    Blue = 8'h61;
end 13'h181d:    begin Red = 8'h4c;    Green = 8'h8f;    Blue = 8'ha9;
end 13'h181e:    begin Red = 8'h48;    Green = 8'h7e;    Blue = 8'h98;
end 13'h181f:    begin Red = 8'h46;    Green = 8'h45;    Blue = 8'h53;
end 13'h1820:    begin Red = 8'h37;    Green = 8'h42;    Blue = 8'h46;
end 13'h1821:    begin Red = 8'h51;    Green = 8'h7f;    Blue = 8'h99;
end 13'h1822:    begin Red = 8'h4e;    Green = 8'h7e;    Blue = 8'h95;
end 13'h1823:    begin Red = 8'h8c;    Green = 8'h6e;    Blue = 8'h25;
end 13'h1824:    begin Red = 8'hc3;    Green = 8'haf;    Blue = 8'h7a;
end 13'h1825:    begin Red = 8'h48;    Green = 8'h2f;    Blue = 8'h42;
end 13'h1826:    begin Red = 8'h2f;    Green = 8'h18;    Blue = 8'h2a;
end 13'h1827:    begin Red = 8'h29;    Green = 8'h18;    Blue = 8'h28;
end 13'h1828:    begin Red = 8'hd2;    Green = 8'hbf;    Blue = 8'h85;
end 13'h1829:    begin Red = 8'haf;    Green = 8'h97;    Blue = 8'h69;
end 13'h182a:    begin Red = 8'h40;    Green = 8'h26;    Blue = 8'h31;
end 13'h182b:    begin Red = 8'h38;    Green = 8'h21;    Blue = 8'h27;
end 13'h182c:    begin Red = 8'h01;    Green = 8'hf1;    Blue = 8'h59;
end 13'h182d:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'h11;
end 13'h182e:    begin Red = 8'h4a;    Green = 8'h28;    Blue = 8'h29;
end 13'h182f:    begin Red = 8'h3e;    Green = 8'h26;    Blue = 8'h34;
end 13'h1830:    begin Red = 8'h38;    Green = 8'h2c;    Blue = 8'h2e;
end 13'h1831:    begin Red = 8'h79;    Green = 8'h48;    Blue = 8'h44;
end 13'h1832:    begin Red = 8'h2d;    Green = 8'h19;    Blue = 8'h1b;
end 13'h1833:    begin Red = 8'h40;    Green = 8'h22;    Blue = 8'h2e;
end 13'h1834:    begin Red = 8'h3c;    Green = 8'h21;    Blue = 8'h26;
end 13'h1835:    begin Red = 8'h33;    Green = 8'h23;    Blue = 8'h24;
end 13'h1836:    begin Red = 8'h33;    Green = 8'h21;    Blue = 8'h21;
end 13'h1837:    begin Red = 8'h00;    Green = 8'h15;    Blue = 8'he8;
end 13'h1838:    begin Red = 8'h63;    Green = 8'h4f;    Blue = 8'h5a;
end 13'h1839:    begin Red = 8'h65;    Green = 8'h58;    Blue = 8'h61;
end 13'h183a:    begin Red = 8'h3b;    Green = 8'h27;    Blue = 8'h28;
end 13'h183b:    begin Red = 8'h00;    Green = 8'h0b;    Blue = 8'h19;
end 13'h183c:    begin Red = 8'hcf;    Green = 8'ha7;    Blue = 8'h21;
end 13'h183d:    begin Red = 8'h2d;    Green = 8'h3c;    Blue = 8'h53;
end 13'h183e:    begin Red = 8'h90;    Green = 8'h9b;    Blue = 8'h8d;
end 13'h183f:    begin Red = 8'hc2;    Green = 8'h64;    Blue = 8'h5a;
end 13'h1840:    begin Red = 8'hc3;    Green = 8'h66;    Blue = 8'h5c;
end 13'h1841:    begin Red = 8'hed;    Green = 8'he0;    Blue = 8'hcb;
end 13'h1842:    begin Red = 8'hbf;    Green = 8'h9e;    Blue = 8'h50;
end 13'h1843:    begin Red = 8'h4c;    Green = 8'h72;    Blue = 8'h84;
end 13'h1844:    begin Red = 8'h54;    Green = 8'h77;    Blue = 8'h8c;
end 13'h1845:    begin Red = 8'h5d;    Green = 8'h58;    Blue = 8'h5d;
end 13'h1846:    begin Red = 8'h75;    Green = 8'hb6;    Blue = 8'hea;
end 13'h1847:    begin Red = 8'h77;    Green = 8'hd1;    Blue = 8'hff;
end 13'h1848:    begin Red = 8'h65;    Green = 8'h55;    Blue = 8'h54;
end 13'h1849:    begin Red = 8'h72;    Green = 8'hbb;    Blue = 8'he6;
end 13'h184a:    begin Red = 8'h5a;    Green = 8'h3f;    Blue = 8'h34;
end 13'h184b:    begin Red = 8'h59;    Green = 8'h43;    Blue = 8'h34;
end 13'h184c:    begin Red = 8'hae;    Green = 8'haf;    Blue = 8'h65;
end 13'h184d:    begin Red = 8'h90;    Green = 8'h84;    Blue = 8'h57;
end 13'h184e:    begin Red = 8'h93;    Green = 8'h88;    Blue = 8'h52;
end 13'h184f:    begin Red = 8'hd9;    Green = 8'hbb;    Blue = 8'h4e;
end 13'h1850:    begin Red = 8'hdd;    Green = 8'hb7;    Blue = 8'h52;
end 13'h1851:    begin Red = 8'hb7;    Green = 8'hbb;    Blue = 8'h92;
end 13'h1852:    begin Red = 8'hb3;    Green = 8'hbb;    Blue = 8'h98;
end 13'h1853:    begin Red = 8'he3;    Green = 8'hc0;    Blue = 8'h88;
end 13'h1854:    begin Red = 8'h00;    Green = 8'h2c;    Blue = 8'he3;
end 13'h1855:    begin Red = 8'h9f;    Green = 8'h9a;    Blue = 8'h63;
end 13'h1856:    begin Red = 8'h93;    Green = 8'h8c;    Blue = 8'h58;
end 13'h1857:    begin Red = 8'h8d;    Green = 8'h87;    Blue = 8'h53;
end 13'h1858:    begin Red = 8'h88;    Green = 8'h85;    Blue = 8'h52;
end 13'h1859:    begin Red = 8'h75;    Green = 8'h76;    Blue = 8'h3d;
end 13'h185a:    begin Red = 8'h68;    Green = 8'h6f;    Blue = 8'h3c;
end 13'h185b:    begin Red = 8'h6e;    Green = 8'h70;    Blue = 8'h3f;
end 13'h185c:    begin Red = 8'h62;    Green = 8'h64;    Blue = 8'h35;
end 13'h185d:    begin Red = 8'h56;    Green = 8'h5e;    Blue = 8'h2d;
end 13'h185e:    begin Red = 8'h59;    Green = 8'h5f;    Blue = 8'h31;
end 13'h185f:    begin Red = 8'hef;    Green = 8'hd6;    Blue = 8'h9e;
end 13'h1860:    begin Red = 8'h04;    Green = 8'h42;    Blue = 8'h90;
end 13'h1861:    begin Red = 8'h8f;    Green = 8'h8c;    Blue = 8'h59;
end 13'h1862:    begin Red = 8'h54;    Green = 8'h52;    Blue = 8'h2c;
end 13'h1863:    begin Red = 8'h49;    Green = 8'h4e;    Blue = 8'h26;
end 13'h1864:    begin Red = 8'h43;    Green = 8'h4f;    Blue = 8'h27;
end 13'h1865:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h99;
end 13'h1866:    begin Red = 8'hc2;    Green = 8'ha1;    Blue = 8'h76;
end 13'h1867:    begin Red = 8'ha9;    Green = 8'h8c;    Blue = 8'h64;
end 13'h1868:    begin Red = 8'h5b;    Green = 8'hc5;    Blue = 8'hc1;
end 13'h1869:    begin Red = 8'h69;    Green = 8'hc9;    Blue = 8'hc7;
end 13'h186a:    begin Red = 8'h29;    Green = 8'h32;    Blue = 8'h43;
end 13'h186b:    begin Red = 8'h4e;    Green = 8'h8a;    Blue = 8'haf;
end 13'h186c:    begin Red = 8'h53;    Green = 8'h91;    Blue = 8'ha6;
end 13'h186d:    begin Red = 8'h2a;    Green = 8'h26;    Blue = 8'h3f;
end 13'h186e:    begin Red = 8'h5a;    Green = 8'h8e;    Blue = 8'hb5;
end 13'h186f:    begin Red = 8'h48;    Green = 8'h79;    Blue = 8'h97;
end 13'h1870:    begin Red = 8'h39;    Green = 8'h75;    Blue = 8'h91;
end 13'h1871:    begin Red = 8'h90;    Green = 8'h65;    Blue = 8'h17;
end 13'h1872:    begin Red = 8'had;    Green = 8'h97;    Blue = 8'h65;
end 13'h1873:    begin Red = 8'hc5;    Green = 8'hb2;    Blue = 8'h78;
end 13'h1874:    begin Red = 8'h4a;    Green = 8'h31;    Blue = 8'h44;
end 13'h1875:    begin Red = 8'h2d;    Green = 8'h19;    Blue = 8'h24;
end 13'h1876:    begin Red = 8'h2c;    Green = 8'h16;    Blue = 8'h23;
end 13'h1877:    begin Red = 8'hd0;    Green = 8'hba;    Blue = 8'h7e;
end 13'h1878:    begin Red = 8'h39;    Green = 8'h29;    Blue = 8'h29;
end 13'h1879:    begin Red = 8'h20;    Green = 8'h15;    Blue = 8'h13;
end 13'h187a:    begin Red = 8'h01;    Green = 8'h81;    Blue = 8'h26;
end 13'h187b:    begin Red = 8'h44;    Green = 8'h2c;    Blue = 8'h2c;
end 13'h187c:    begin Red = 8'h36;    Green = 8'h25;    Blue = 8'h2d;
end 13'h187d:    begin Red = 8'h7b;    Green = 8'h47;    Blue = 8'h4b;
end 13'h187e:    begin Red = 8'h5e;    Green = 8'h52;    Blue = 8'h5e;
end 13'h187f:    begin Red = 8'h5c;    Green = 8'h4f;    Blue = 8'h56;
end 13'h1880:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h38;
end 13'h1881:    begin Red = 8'h00;    Green = 8'h1a;    Blue = 8'hd7;
end 13'h1882:    begin Red = 8'h67;    Green = 8'h5a;    Blue = 8'h64;
end 13'h1883:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'h5a;
end 13'h1884:    begin Red = 8'hfc;    Green = 8'hc3;    Blue = 8'h2b;
end 13'h1885:    begin Red = 8'h42;    Green = 8'h43;    Blue = 8'h58;
end 13'h1886:    begin Red = 8'hd2;    Green = 8'h64;    Blue = 8'h5c;
end 13'h1887:    begin Red = 8'hd4;    Green = 8'h61;    Blue = 8'h5e;
end 13'h1888:    begin Red = 8'hd4;    Green = 8'h63;    Blue = 8'h5a;
end 13'h1889:    begin Red = 8'hbe;    Green = 8'h4b;    Blue = 8'h44;
end 13'h188a:    begin Red = 8'hba;    Green = 8'ha7;    Blue = 8'h5a;
end 13'h188b:    begin Red = 8'h5d;    Green = 8'h71;    Blue = 8'h91;
end 13'h188c:    begin Red = 8'h55;    Green = 8'h80;    Blue = 8'h98;
end 13'h188d:    begin Red = 8'h5a;    Green = 8'h7f;    Blue = 8'h95;
end 13'h188e:    begin Red = 8'h75;    Green = 8'hc3;    Blue = 8'hf7;
end 13'h188f:    begin Red = 8'h71;    Green = 8'hc3;    Blue = 8'hf2;
end 13'h1890:    begin Red = 8'h6e;    Green = 8'h57;    Blue = 8'h51;
end 13'h1891:    begin Red = 8'h63;    Green = 8'h45;    Blue = 8'h3e;
end 13'h1892:    begin Red = 8'h75;    Green = 8'hbb;    Blue = 8'hf6;
end 13'h1893:    begin Red = 8'hac;    Green = 8'hb1;    Blue = 8'h50;
end 13'h1894:    begin Red = 8'hbb;    Green = 8'hbe;    Blue = 8'h65;
end 13'h1895:    begin Red = 8'h74;    Green = 8'h71;    Blue = 8'h4e;
end 13'h1896:    begin Red = 8'hf5;    Green = 8'hca;    Blue = 8'h50;
end 13'h1897:    begin Red = 8'hfa;    Green = 8'hce;    Blue = 8'h52;
end 13'h1898:    begin Red = 8'h5f;    Green = 8'h60;    Blue = 8'h64;
end 13'h1899:    begin Red = 8'h8c;    Green = 8'h88;    Blue = 8'h73;
end 13'h189a:    begin Red = 8'hf7;    Green = 8'hd7;    Blue = 8'ha4;
end 13'h189b:    begin Red = 8'hf2;    Green = 8'hd2;    Blue = 8'h9f;
end 13'h189c:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h21;
end 13'h189d:    begin Red = 8'h04;    Green = 8'ha2;    Blue = 8'he0;
end 13'h189e:    begin Red = 8'h9b;    Green = 8'h94;    Blue = 8'h5e;
end 13'h189f:    begin Red = 8'h8d;    Green = 8'h89;    Blue = 8'h59;
end 13'h18a0:    begin Red = 8'h71;    Green = 8'h71;    Blue = 8'h3d;
end 13'h18a1:    begin Red = 8'h6d;    Green = 8'h65;    Blue = 8'h36;
end 13'h18a2:    begin Red = 8'h5f;    Green = 8'h5e;    Blue = 8'h2e;
end 13'h18a3:    begin Red = 8'h5e;    Green = 8'h62;    Blue = 8'h30;
end 13'h18a4:    begin Red = 8'h06;    Green = 8'h84;    Blue = 8'h24;
end 13'h18a5:    begin Red = 8'hfa;    Green = 8'he0;    Blue = 8'ha5;
end 13'h18a6:    begin Red = 8'he0;    Green = 8'hbf;    Blue = 8'h8a;
end 13'h18a7:    begin Red = 8'he5;    Green = 8'hca;    Blue = 8'h95;
end 13'h18a8:    begin Red = 8'hdd;    Green = 8'hb7;    Blue = 8'h86;
end 13'h18a9:    begin Red = 8'hde;    Green = 8'hbe;    Blue = 8'h83;
end 13'h18aa:    begin Red = 8'hc0;    Green = 8'ha0;    Blue = 8'h6d;
end 13'h18ab:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'hb6;
end 13'h18ac:    begin Red = 8'h61;    Green = 8'h5e;    Blue = 8'h3b;
end 13'h18ad:    begin Red = 8'hd1;    Green = 8'hdb;    Blue = 8'hb7;
end 13'h18ae:    begin Red = 8'h60;    Green = 8'h61;    Blue = 8'h35;
end 13'h18af:    begin Red = 8'hb3;    Green = 8'h98;    Blue = 8'h6b;
end 13'h18b0:    begin Red = 8'h35;    Green = 8'h34;    Blue = 8'h39;
end 13'h18b1:    begin Red = 8'he7;    Green = 8'hec;    Blue = 8'he8;
end 13'h18b2:    begin Red = 8'h85;    Green = 8'hd0;    Blue = 8'hd6;
end 13'h18b3:    begin Red = 8'h2a;    Green = 8'h35;    Blue = 8'h3b;
end 13'h18b4:    begin Red = 8'h39;    Green = 8'h4f;    Blue = 8'h5d;
end 13'h18b5:    begin Red = 8'h95;    Green = 8'heb;    Blue = 8'hea;
end 13'h18b6:    begin Red = 8'h96;    Green = 8'he7;    Blue = 8'hea;
end 13'h18b7:    begin Red = 8'h41;    Green = 8'h4c;    Blue = 8'h60;
end 13'h18b8:    begin Red = 8'h95;    Green = 8'hea;    Blue = 8'hef;
end 13'h18b9:    begin Red = 8'h80;    Green = 8'hce;    Blue = 8'hd2;
end 13'h18ba:    begin Red = 8'hc7;    Green = 8'hb2;    Blue = 8'h7b;
end 13'h18bb:    begin Red = 8'h32;    Green = 8'h1e;    Blue = 8'h2a;
end 13'h18bc:    begin Red = 8'h2f;    Green = 8'h1e;    Blue = 8'h28;
end 13'h18bd:    begin Red = 8'h31;    Green = 8'h1c;    Blue = 8'h2d;
end 13'h18be:    begin Red = 8'hcb;    Green = 8'hb7;    Blue = 8'h7c;
end 13'h18bf:    begin Red = 8'h3a;    Green = 8'h23;    Blue = 8'h29;
end 13'h18c0:    begin Red = 8'h3a;    Green = 8'h25;    Blue = 8'h2c;
end 13'h18c1:    begin Red = 8'h7a;    Green = 8'h46;    Blue = 8'h48;
end 13'h18c2:    begin Red = 8'h2a;    Green = 8'h1f;    Blue = 8'h25;
end 13'h18c3:    begin Red = 8'h77;    Green = 8'h42;    Blue = 8'h4a;
end 13'h18c4:    begin Red = 8'h53;    Green = 8'h4c;    Blue = 8'h53;
end 13'h18c5:    begin Red = 8'h59;    Green = 8'h4d;    Blue = 8'h59;
end 13'h18c6:    begin Red = 8'h41;    Green = 8'h2a;    Blue = 8'h32;
end 13'h18c7:    begin Red = 8'h63;    Green = 8'h56;    Blue = 8'h5d;
end 13'h18c8:    begin Red = 8'h3d;    Green = 8'h24;    Blue = 8'h2a;
end 13'h18c9:    begin Red = 8'h36;    Green = 8'h20;    Blue = 8'h23;
end 13'h18ca:    begin Red = 8'h00;    Green = 8'h0f;    Blue = 8'h2c;
end 13'h18cb:    begin Red = 8'h2e;    Green = 8'h2e;    Blue = 8'h2e;
end 13'h18cc:    begin Red = 8'h27;    Green = 8'h25;    Blue = 8'h28;
end 13'h18cd:    begin Red = 8'hd0;    Green = 8'ha8;    Blue = 8'h25;
end 13'h18ce:    begin Red = 8'h4d;    Green = 8'h4f;    Blue = 8'h4e;
end 13'h18cf:    begin Red = 8'haa;    Green = 8'ha3;    Blue = 8'h9f;
end 13'h18d0:    begin Red = 8'h5d;    Green = 8'h58;    Blue = 8'h4a;
end 13'h18d1:    begin Red = 8'h67;    Green = 8'h88;    Blue = 8'h9e;
end 13'h18d2:    begin Red = 8'h6d;    Green = 8'h98;    Blue = 8'hb5;
end 13'h18d3:    begin Red = 8'h4e;    Green = 8'h4b;    Blue = 8'h42;
end 13'h18d4:    begin Red = 8'h68;    Green = 8'h8b;    Blue = 8'ha2;
end 13'h18d5:    begin Red = 8'h67;    Green = 8'h87;    Blue = 8'ha3;
end 13'h18d6:    begin Red = 8'h6c;    Green = 8'hb7;    Blue = 8'he7;
end 13'h18d7:    begin Red = 8'ha0;    Green = 8'h89;    Blue = 8'h55;
end 13'h18d8:    begin Red = 8'hea;    Green = 8'he1;    Blue = 8'hcf;
end 13'h18d9:    begin Red = 8'h78;    Green = 8'h79;    Blue = 8'h75;
end 13'h18da:    begin Red = 8'hd7;    Green = 8'hba;    Blue = 8'h52;
end 13'h18db:    begin Red = 8'h3d;    Green = 8'h3b;    Blue = 8'h4e;
end 13'h18dc:    begin Red = 8'h76;    Green = 8'h72;    Blue = 8'h70;
end 13'h18dd:    begin Red = 8'h73;    Green = 8'h73;    Blue = 8'h79;
end 13'h18de:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'hd0;
end 13'h18df:    begin Red = 8'h6b;    Green = 8'h6c;    Blue = 8'h40;
end 13'h18e0:    begin Red = 8'h5e;    Green = 8'h5c;    Blue = 8'h35;
end 13'h18e1:    begin Red = 8'h51;    Green = 8'h57;    Blue = 8'h29;
end 13'h18e2:    begin Red = 8'h52;    Green = 8'h50;    Blue = 8'h29;
end 13'h18e3:    begin Red = 8'h50;    Green = 8'h52;    Blue = 8'h2a;
end 13'h18e4:    begin Red = 8'h06;    Green = 8'h33;    Blue = 8'hf5;
end 13'h18e5:    begin Red = 8'h04;    Green = 8'h02;    Blue = 8'h90;
end 13'h18e6:    begin Red = 8'h4f;    Green = 8'h50;    Blue = 8'h2e;
end 13'h18e7:    begin Red = 8'h46;    Green = 8'h47;    Blue = 8'h25;
end 13'h18e8:    begin Red = 8'h42;    Green = 8'h43;    Blue = 8'h24;
end 13'h18e9:    begin Red = 8'h3f;    Green = 8'h43;    Blue = 8'h22;
end 13'h18ea:    begin Red = 8'h05;    Green = 8'h33;    Blue = 8'h45;
end 13'h18eb:    begin Red = 8'h54;    Green = 8'h55;    Blue = 8'h5a;
end 13'h18ec:    begin Red = 8'hb8;    Green = 8'hdb;    Blue = 8'hd5;
end 13'h18ed:    begin Red = 8'h7a;    Green = 8'hc7;    Blue = 8'hd7;
end 13'h18ee:    begin Red = 8'h8c;    Green = 8'hcb;    Blue = 8'hd0;
end 13'h18ef:    begin Red = 8'h82;    Green = 8'hcc;    Blue = 8'hcf;
end 13'h18f0:    begin Red = 8'h81;    Green = 8'hcf;    Blue = 8'hd9;
end 13'h18f1:    begin Red = 8'h86;    Green = 8'hcd;    Blue = 8'hd3;
end 13'h18f2:    begin Red = 8'h36;    Green = 8'h21;    Blue = 8'h32;
end 13'h18f3:    begin Red = 8'h37;    Green = 8'h22;    Blue = 8'h35;
end 13'h18f4:    begin Red = 8'h48;    Green = 8'h2e;    Blue = 8'h39;
end 13'h18f5:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'h2e;
end 13'h18f6:    begin Red = 8'h00;    Green = 8'h12;    Blue = 8'hb1;
end 13'h18f7:    begin Red = 8'h4a;    Green = 8'h30;    Blue = 8'h3d;
end 13'h18f8:    begin Red = 8'h4a;    Green = 8'h2a;    Blue = 8'h39;
end 13'h18f9:    begin Red = 8'h42;    Green = 8'h2e;    Blue = 8'h39;
end 13'h18fa:    begin Red = 8'h3d;    Green = 8'h2d;    Blue = 8'h38;
end 13'h18fb:    begin Red = 8'h41;    Green = 8'h22;    Blue = 8'h32;
end 13'h18fc:    begin Red = 8'h35;    Green = 8'h25;    Blue = 8'h32;
end 13'h18fd:    begin Red = 8'h3b;    Green = 8'h29;    Blue = 8'h35;
end 13'h18fe:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'h3a;
end 13'h18ff:    begin Red = 8'h50;    Green = 8'h34;    Blue = 8'h42;
end 13'h1900:    begin Red = 8'h44;    Green = 8'h30;    Blue = 8'h3b;
end 13'h1901:    begin Red = 8'h3f;    Green = 8'h29;    Blue = 8'h36;
end 13'h1902:    begin Red = 8'h01;    Green = 8'h23;    Blue = 8'h16;
end 13'h1903:    begin Red = 8'hf0;    Green = 8'hd3;    Blue = 8'hb1;
end 13'h1904:    begin Red = 8'h56;    Green = 8'h4b;    Blue = 8'h45;
end 13'h1905:    begin Red = 8'h70;    Green = 8'hb7;    Blue = 8'he6;
end 13'h1906:    begin Red = 8'h78;    Green = 8'hc7;    Blue = 8'hfd;
end 13'h1907:    begin Red = 8'h55;    Green = 8'h75;    Blue = 8'h89;
end 13'h1908:    begin Red = 8'h63;    Green = 8'h87;    Blue = 8'ha1;
end 13'h1909:    begin Red = 8'h61;    Green = 8'h8d;    Blue = 8'h99;
end 13'h190a:    begin Red = 8'h61;    Green = 8'h85;    Blue = 8'h9a;
end 13'h190b:    begin Red = 8'h64;    Green = 8'h87;    Blue = 8'h9b;
end 13'h190c:    begin Red = 8'h62;    Green = 8'h8c;    Blue = 8'ha7;
end 13'h190d:    begin Red = 8'hfc;    Green = 8'h70;    Blue = 8'h4f;
end 13'h190e:    begin Red = 8'hf4;    Green = 8'h78;    Blue = 8'h64;
end 13'h190f:    begin Red = 8'h75;    Green = 8'h74;    Blue = 8'h53;
end 13'h1910:    begin Red = 8'h78;    Green = 8'h70;    Blue = 8'h6f;
end 13'h1911:    begin Red = 8'h6f;    Green = 8'h71;    Blue = 8'h6c;
end 13'h1912:    begin Red = 8'h77;    Green = 8'h75;    Blue = 8'h71;
end 13'h1913:    begin Red = 8'h04;    Green = 8'hf2;    Blue = 8'he1;
end 13'h1914:    begin Red = 8'h68;    Green = 8'h65;    Blue = 8'h38;
end 13'h1915:    begin Red = 8'h5b;    Green = 8'h5e;    Blue = 8'h2f;
end 13'h1916:    begin Red = 8'h59;    Green = 8'h58;    Blue = 8'h2a;
end 13'h1917:    begin Red = 8'h58;    Green = 8'h5b;    Blue = 8'h2e;
end 13'h1918:    begin Red = 8'h06;    Green = 8'h54;    Blue = 8'h09;
end 13'h1919:    begin Red = 8'hea;    Green = 8'hb9;    Blue = 8'h7e;
end 13'h191a:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'hc3;
end 13'h191b:    begin Red = 8'h5d;    Green = 8'h5a;    Blue = 8'h37;
end 13'h191c:    begin Red = 8'h8a;    Green = 8'h83;    Blue = 8'h55;
end 13'h191d:    begin Red = 8'h84;    Green = 8'h7e;    Blue = 8'h4e;
end 13'h191e:    begin Red = 8'h75;    Green = 8'h70;    Blue = 8'h4a;
end 13'h191f:    begin Red = 8'h48;    Green = 8'h4a;    Blue = 8'h22;
end 13'h1920:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h57;
end 13'h1921:    begin Red = 8'h48;    Green = 8'h40;    Blue = 8'h4b;
end 13'h1922:    begin Red = 8'h36;    Green = 8'h31;    Blue = 8'h38;
end 13'h1923:    begin Red = 8'hb5;    Green = 8'hdd;    Blue = 8'hd5;
end 13'h1924:    begin Red = 8'h6e;    Green = 8'hcd;    Blue = 8'hc7;
end 13'h1925:    begin Red = 8'h79;    Green = 8'hca;    Blue = 8'hcd;
end 13'h1926:    begin Red = 8'h74;    Green = 8'hd1;    Blue = 8'hd9;
end 13'h1927:    begin Red = 8'h73;    Green = 8'he6;    Blue = 8'hed;
end 13'h1928:    begin Red = 8'h76;    Green = 8'he3;    Blue = 8'hea;
end 13'h1929:    begin Red = 8'h74;    Green = 8'he9;    Blue = 8'hf3;
end 13'h192a:    begin Red = 8'h07;    Green = 8'hf6;    Blue = 8'hdb;
end 13'h192b:    begin Red = 8'h08;    Green = 8'h66;    Blue = 8'h37;
end 13'h192c:    begin Red = 8'h4d;    Green = 8'h30;    Blue = 8'h46;
end 13'h192d:    begin Red = 8'h35;    Green = 8'h22;    Blue = 8'h26;
end 13'h192e:    begin Red = 8'h33;    Green = 8'h21;    Blue = 8'h2d;
end 13'h192f:    begin Red = 8'h35;    Green = 8'h1f;    Blue = 8'h2b;
end 13'h1930:    begin Red = 8'h34;    Green = 8'h1e;    Blue = 8'h35;
end 13'h1931:    begin Red = 8'hf3;    Green = 8'hff;    Blue = 8'hca;
end 13'h1932:    begin Red = 8'h46;    Green = 8'h32;    Blue = 8'h31;
end 13'h1933:    begin Red = 8'h35;    Green = 8'h14;    Blue = 8'h25;
end 13'h1934:    begin Red = 8'h29;    Green = 8'h12;    Blue = 8'h1a;
end 13'h1935:    begin Red = 8'h42;    Green = 8'h2d;    Blue = 8'h34;
end 13'h1936:    begin Red = 8'h01;    Green = 8'h81;    Blue = 8'h30;
end 13'h1937:    begin Red = 8'h51;    Green = 8'h36;    Blue = 8'h3b;
end 13'h1938:    begin Red = 8'h47;    Green = 8'h32;    Blue = 8'h39;
end 13'h1939:    begin Red = 8'h01;    Green = 8'h36;    Blue = 8'h17;
end 13'h193a:    begin Red = 8'h34;    Green = 8'h33;    Blue = 8'h31;
end 13'h193b:    begin Red = 8'h35;    Green = 8'h38;    Blue = 8'h3d;
end 13'h193c:    begin Red = 8'h4a;    Green = 8'h4a;    Blue = 8'h4a;
end 13'h193d:    begin Red = 8'h31;    Green = 8'h36;    Blue = 8'h3c;
end 13'h193e:    begin Red = 8'hfc;    Green = 8'hf2;    Blue = 8'hb7;
end 13'h193f:    begin Red = 8'h7d;    Green = 8'hc8;    Blue = 8'hfb;
end 13'h1940:    begin Red = 8'h7d;    Green = 8'hd2;    Blue = 8'hff;
end 13'h1941:    begin Red = 8'h59;    Green = 8'h75;    Blue = 8'h84;
end 13'h1942:    begin Red = 8'h55;    Green = 8'h71;    Blue = 8'h80;
end 13'h1943:    begin Red = 8'h4f;    Green = 8'h78;    Blue = 8'h83;
end 13'h1944:    begin Red = 8'h5d;    Green = 8'h78;    Blue = 8'h8f;
end 13'h1945:    begin Red = 8'h4b;    Green = 8'h69;    Blue = 8'h78;
end 13'h1946:    begin Red = 8'h52;    Green = 8'h70;    Blue = 8'h85;
end 13'h1947:    begin Red = 8'h6b;    Green = 8'h8c;    Blue = 8'ha0;
end 13'h1948:    begin Red = 8'h64;    Green = 8'h84;    Blue = 8'h9e;
end 13'h1949:    begin Red = 8'h62;    Green = 8'h89;    Blue = 8'ha3;
end 13'h194a:    begin Red = 8'h6b;    Green = 8'h93;    Blue = 8'haf;
end 13'h194b:    begin Red = 8'h6c;    Green = 8'h96;    Blue = 8'hb9;
end 13'h194c:    begin Red = 8'h68;    Green = 8'h84;    Blue = 8'h9d;
end 13'h194d:    begin Red = 8'h5e;    Green = 8'h8c;    Blue = 8'ha1;
end 13'h194e:    begin Red = 8'h63;    Green = 8'h8c;    Blue = 8'h9e;
end 13'h194f:    begin Red = 8'h47;    Green = 8'h8f;    Blue = 8'hac;
end 13'h1950:    begin Red = 8'hff;    Green = 8'h61;    Blue = 8'h49;
end 13'h1951:    begin Red = 8'hfa;    Green = 8'h5b;    Blue = 8'h4f;
end 13'h1952:    begin Red = 8'hbe;    Green = 8'hc2;    Blue = 8'h6a;
end 13'h1953:    begin Red = 8'he9;    Green = 8'hd9;    Blue = 8'hc5;
end 13'h1954:    begin Red = 8'h59;    Green = 8'h5a;    Blue = 8'h5b;
end 13'h1955:    begin Red = 8'h62;    Green = 8'h61;    Blue = 8'h69;
end 13'h1956:    begin Red = 8'h03;    Green = 8'h01;    Blue = 8'h40;
end 13'h1957:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'hc4;
end 13'h1958:    begin Red = 8'h95;    Green = 8'h8e;    Blue = 8'h5a;
end 13'h1959:    begin Red = 8'h70;    Green = 8'h6f;    Blue = 8'h41;
end 13'h195a:    begin Red = 8'h59;    Green = 8'h60;    Blue = 8'h2d;
end 13'h195b:    begin Red = 8'h5b;    Green = 8'h5a;    Blue = 8'h2c;
end 13'h195c:    begin Red = 8'h6a;    Green = 8'h5a;    Blue = 8'h36;
end 13'h195d:    begin Red = 8'h56;    Green = 8'h56;    Blue = 8'h30;
end 13'h195e:    begin Red = 8'h4b;    Green = 8'h4b;    Blue = 8'h27;
end 13'h195f:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h45;
end 13'h1960:    begin Red = 8'h8c;    Green = 8'h94;    Blue = 8'h7d;
end 13'h1961:    begin Red = 8'he2;    Green = 8'he2;    Blue = 8'hea;
end 13'h1962:    begin Red = 8'hb7;    Green = 8'hda;    Blue = 8'hde;
end 13'h1963:    begin Red = 8'hb4;    Green = 8'hde;    Blue = 8'hd0;
end 13'h1964:    begin Red = 8'hbb;    Green = 8'hd9;    Blue = 8'he1;
end 13'h1965:    begin Red = 8'hbe;    Green = 8'he1;    Blue = 8'he5;
end 13'h1966:    begin Red = 8'hb2;    Green = 8'hf2;    Blue = 8'hfb;
end 13'h1967:    begin Red = 8'hbd;    Green = 8'h64;    Blue = 8'h66;
end 13'h1968:    begin Red = 8'hbd;    Green = 8'h62;    Blue = 8'h61;
end 13'h1969:    begin Red = 8'hc1;    Green = 8'h67;    Blue = 8'h69;
end 13'h196a:    begin Red = 8'h08;    Green = 8'h46;    Blue = 8'h15;
end 13'h196b:    begin Red = 8'h3c;    Green = 8'h27;    Blue = 8'h2e;
end 13'h196c:    begin Red = 8'h3d;    Green = 8'h28;    Blue = 8'h31;
end 13'h196d:    begin Red = 8'h3d;    Green = 8'h25;    Blue = 8'h3b;
end 13'h196e:    begin Red = 8'hca;    Green = 8'hb4;    Blue = 8'h7b;
end 13'h196f:    begin Red = 8'h73;    Green = 8'h65;    Blue = 8'h4b;
end 13'h1970:    begin Red = 8'hfb;    Green = 8'hf7;    Blue = 8'hba;
end 13'h1971:    begin Red = 8'h57;    Green = 8'h2c;    Blue = 8'h47;
end 13'h1972:    begin Red = 8'hea;    Green = 8'hf5;    Blue = 8'hc4;
end 13'h1973:    begin Red = 8'h3e;    Green = 8'h22;    Blue = 8'h39;
end 13'h1974:    begin Red = 8'h3b;    Green = 8'h23;    Blue = 8'h33;
end 13'h1975:    begin Red = 8'h3a;    Green = 8'h24;    Blue = 8'h39;
end 13'h1976:    begin Red = 8'h02;    Green = 8'h01;    Blue = 8'h5f;
end 13'h1977:    begin Red = 8'h48;    Green = 8'h2a;    Blue = 8'h42;
end 13'h1978:    begin Red = 8'h45;    Green = 8'h27;    Blue = 8'h3f;
end 13'h1979:    begin Red = 8'h41;    Green = 8'h25;    Blue = 8'h3c;
end 13'h197a:    begin Red = 8'h3c;    Green = 8'h25;    Blue = 8'h37;
end 13'h197b:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h02;
end 13'h197c:    begin Red = 8'h42;    Green = 8'h27;    Blue = 8'h38;
end 13'h197d:    begin Red = 8'h3f;    Green = 8'h26;    Blue = 8'h39;
end 13'h197e:    begin Red = 8'h00;    Green = 8'he2;    Blue = 8'h18;
end 13'h197f:    begin Red = 8'hfd;    Green = 8'hf1;    Blue = 8'hc1;
end 13'h1980:    begin Red = 8'h73;    Green = 8'h66;    Blue = 8'h67;
end 13'h1981:    begin Red = 8'h7b;    Green = 8'h74;    Blue = 8'h6e;
end 13'h1982:    begin Red = 8'h88;    Green = 8'h85;    Blue = 8'h6e;
end 13'h1983:    begin Red = 8'hd2;    Green = 8'hcd;    Blue = 8'hbe;
end 13'h1984:    begin Red = 8'h50;    Green = 8'h74;    Blue = 8'h86;
end 13'h1985:    begin Red = 8'h52;    Green = 8'h75;    Blue = 8'h78;
end 13'h1986:    begin Red = 8'h7d;    Green = 8'hbf;    Blue = 8'hfd;
end 13'h1987:    begin Red = 8'h60;    Green = 8'h7d;    Blue = 8'h84;
end 13'h1988:    begin Red = 8'h4a;    Green = 8'h90;    Blue = 8'haf;
end 13'h1989:    begin Red = 8'hee;    Green = 8'h71;    Blue = 8'h64;
end 13'h198a:    begin Red = 8'he0;    Green = 8'hf7;    Blue = 8'hde;
end 13'h198b:    begin Red = 8'h9a;    Green = 8'h8b;    Blue = 8'h5c;
end 13'h198c:    begin Red = 8'h04;    Green = 8'ha2;    Blue = 8'hd5;
end 13'h198d:    begin Red = 8'h9d;    Green = 8'h96;    Blue = 8'h5f;
end 13'h198e:    begin Red = 8'h7c;    Green = 8'h79;    Blue = 8'h44;
end 13'h198f:    begin Red = 8'h79;    Green = 8'h72;    Blue = 8'h44;
end 13'h1990:    begin Red = 8'h69;    Green = 8'h6a;    Blue = 8'h3e;
end 13'h1991:    begin Red = 8'h55;    Green = 8'h58;    Blue = 8'h2b;
end 13'h1992:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'h91;
end 13'h1993:    begin Red = 8'h6b;    Green = 8'h63;    Blue = 8'h34;
end 13'h1994:    begin Red = 8'hce;    Green = 8'hd7;    Blue = 8'hb5;
end 13'h1995:    begin Red = 8'h53;    Green = 8'h54;    Blue = 8'h32;
end 13'h1996:    begin Red = 8'h05;    Green = 8'h23;    Blue = 8'h34;
end 13'h1997:    begin Red = 8'h87;    Green = 8'h67;    Blue = 8'h14;
end 13'h1998:    begin Red = 8'h8a;    Green = 8'h8e;    Blue = 8'h9a;
end 13'h1999:    begin Red = 8'heb;    Green = 8'hf3;    Blue = 8'hf6;
end 13'h199a:    begin Red = 8'hb3;    Green = 8'hd8;    Blue = 8'hd1;
end 13'h199b:    begin Red = 8'hb6;    Green = 8'hde;    Blue = 8'hde;
end 13'h199c:    begin Red = 8'hc1;    Green = 8'h37;    Blue = 8'h2a;
end 13'h199d:    begin Red = 8'hbd;    Green = 8'h4c;    Blue = 8'h48;
end 13'h199e:    begin Red = 8'hbb;    Green = 8'h62;    Blue = 8'h5e;
end 13'h199f:    begin Red = 8'hbe;    Green = 8'h61;    Blue = 8'h5a;
end 13'h19a0:    begin Red = 8'hb6;    Green = 8'h64;    Blue = 8'h59;
end 13'h19a1:    begin Red = 8'h88;    Green = 8'h69;    Blue = 8'h19;
end 13'h19a2:    begin Red = 8'hff;    Green = 8'hf4;    Blue = 8'hbc;
end 13'h19a3:    begin Red = 8'h4c;    Green = 8'h2d;    Blue = 8'h56;
end 13'h19a4:    begin Red = 8'he7;    Green = 8'hf6;    Blue = 8'hc2;
end 13'h19a5:    begin Red = 8'h3e;    Green = 8'h23;    Blue = 8'h44;
end 13'h19a6:    begin Red = 8'h3b;    Green = 8'h1e;    Blue = 8'h3d;
end 13'h19a7:    begin Red = 8'h01;    Green = 8'hd1;    Blue = 8'h4b;
end 13'h19a8:    begin Red = 8'h00;    Green = 8'h16;    Blue = 8'hf5;
end 13'h19a9:    begin Red = 8'h4b;    Green = 8'h2b;    Blue = 8'h50;
end 13'h19aa:    begin Red = 8'h49;    Green = 8'h2b;    Blue = 8'h4d;
end 13'h19ab:    begin Red = 8'h46;    Green = 8'h29;    Blue = 8'h48;
end 13'h19ac:    begin Red = 8'h40;    Green = 8'h27;    Blue = 8'h45;
end 13'h19ad:    begin Red = 8'h40;    Green = 8'h25;    Blue = 8'h48;
end 13'h19ae:    begin Red = 8'h3c;    Green = 8'h23;    Blue = 8'h41;
end 13'h19af:    begin Red = 8'h3a;    Green = 8'h1f;    Blue = 8'h40;
end 13'h19b0:    begin Red = 8'h46;    Green = 8'h26;    Blue = 8'h4b;
end 13'h19b1:    begin Red = 8'h42;    Green = 8'h29;    Blue = 8'h47;
end 13'h19b2:    begin Red = 8'h00;    Green = 8'he0;    Blue = 8'h1e;
end 13'h19b3:    begin Red = 8'hd6;    Green = 8'hb8;    Blue = 8'h82;
end 13'h19b4:    begin Red = 8'h8c;    Green = 8'h8d;    Blue = 8'h89;
end 13'h19b5:    begin Red = 8'h63;    Green = 8'h61;    Blue = 8'h5b;
end 13'h19b6:    begin Red = 8'hc5;    Green = 8'haf;    Blue = 8'h83;
end 13'h19b7:    begin Red = 8'h88;    Green = 8'h78;    Blue = 8'h70;
end 13'h19b8:    begin Red = 8'h83;    Green = 8'h86;    Blue = 8'h5e;
end 13'h19b9:    begin Red = 8'hd2;    Green = 8'hb8;    Blue = 8'h7b;
end 13'h19ba:    begin Red = 8'hd6;    Green = 8'hb7;    Blue = 8'h7d;
end 13'h19bb:    begin Red = 8'h61;    Green = 8'h71;    Blue = 8'h87;
end 13'h19bc:    begin Red = 8'h53;    Green = 8'h78;    Blue = 8'h92;
end 13'h19bd:    begin Red = 8'h64;    Green = 8'h8e;    Blue = 8'ha9;
end 13'h19be:    begin Red = 8'h62;    Green = 8'h88;    Blue = 8'h9e;
end 13'h19bf:    begin Red = 8'haf;    Green = 8'hb9;    Blue = 8'hbe;
end 13'h19c0:    begin Red = 8'hb4;    Green = 8'hb8;    Blue = 8'hbd;
end 13'h19c1:    begin Red = 8'haf;    Green = 8'hbb;    Blue = 8'hbb;
end 13'h19c2:    begin Red = 8'ha7;    Green = 8'hab;    Blue = 8'hb2;
end 13'h19c3:    begin Red = 8'h79;    Green = 8'hcd;    Blue = 8'hfb;
end 13'h19c4:    begin Red = 8'h78;    Green = 8'hc1;    Blue = 8'hfd;
end 13'h19c5:    begin Red = 8'h64;    Green = 8'h80;    Blue = 8'h91;
end 13'h19c6:    begin Red = 8'h47;    Green = 8'h80;    Blue = 8'haf;
end 13'h19c7:    begin Red = 8'hb9;    Green = 8'hd7;    Blue = 8'h54;
end 13'h19c8:    begin Red = 8'he7;    Green = 8'hec;    Blue = 8'he1;
end 13'h19c9:    begin Red = 8'hc3;    Green = 8'hcd;    Blue = 8'hbb;
end 13'h19ca:    begin Red = 8'hcc;    Green = 8'hc8;    Blue = 8'hb9;
end 13'h19cb:    begin Red = 8'hca;    Green = 8'hca;    Blue = 8'hb2;
end 13'h19cc:    begin Red = 8'h04;    Green = 8'h62;    Blue = 8'hd4;
end 13'h19cd:    begin Red = 8'h77;    Green = 8'h74;    Blue = 8'h41;
end 13'h19ce:    begin Red = 8'h5f;    Green = 8'h67;    Blue = 8'h36;
end 13'h19cf:    begin Red = 8'h68;    Green = 8'h61;    Blue = 8'h35;
end 13'h19d0:    begin Red = 8'h53;    Green = 8'h5b;    Blue = 8'h2c;
end 13'h19d1:    begin Red = 8'h06;    Green = 8'h43;    Blue = 8'hf8;
end 13'h19d2:    begin Red = 8'h83;    Green = 8'h82;    Blue = 8'h4c;
end 13'h19d3:    begin Red = 8'h66;    Green = 8'h60;    Blue = 8'h30;
end 13'h19d4:    begin Red = 8'h4d;    Green = 8'h4f;    Blue = 8'h27;
end 13'h19d5:    begin Red = 8'h44;    Green = 8'h4a;    Blue = 8'h24;
end 13'h19d6:    begin Red = 8'hcf;    Green = 8'hd4;    Blue = 8'haf;
end 13'h19d7:    begin Red = 8'h82;    Green = 8'h93;    Blue = 8'h9a;
end 13'h19d8:    begin Red = 8'h7c;    Green = 8'h90;    Blue = 8'h97;
end 13'h19d9:    begin Red = 8'he0;    Green = 8'he6;    Blue = 8'he6;
end 13'h19da:    begin Red = 8'hae;    Green = 8'hd7;    Blue = 8'hdb;
end 13'h19db:    begin Red = 8'hb8;    Green = 8'hd7;    Blue = 8'hda;
end 13'h19dc:    begin Red = 8'hbb;    Green = 8'h4a;    Blue = 8'h3a;
end 13'h19dd:    begin Red = 8'hc4;    Green = 8'h62;    Blue = 8'h55;
end 13'h19de:    begin Red = 8'hf1;    Green = 8'hd0;    Blue = 8'had;
end 13'h19df:    begin Red = 8'h44;    Green = 8'h2f;    Blue = 8'h2e;
end 13'h19e0:    begin Red = 8'h40;    Green = 8'h2f;    Blue = 8'h37;
end 13'h19e1:    begin Red = 8'h42;    Green = 8'h2a;    Blue = 8'h42;
end 13'h19e2:    begin Red = 8'h41;    Green = 8'h29;    Blue = 8'h3f;
end 13'h19e3:    begin Red = 8'hfd;    Green = 8'hfa;    Blue = 8'hb7;
end 13'h19e4:    begin Red = 8'h4b;    Green = 8'h30;    Blue = 8'h51;
end 13'h19e5:    begin Red = 8'he5;    Green = 8'hf3;    Blue = 8'hc2;
end 13'h19e6:    begin Red = 8'h3d;    Green = 8'h21;    Blue = 8'h47;
end 13'h19e7:    begin Red = 8'h48;    Green = 8'h2d;    Blue = 8'h3e;
end 13'h19e8:    begin Red = 8'h46;    Green = 8'h2d;    Blue = 8'h4b;
end 13'h19e9:    begin Red = 8'h42;    Green = 8'h25;    Blue = 8'h43;
end 13'h19ea:    begin Red = 8'h3a;    Green = 8'h27;    Blue = 8'h3d;
end 13'h19eb:    begin Red = 8'h35;    Green = 8'h1c;    Blue = 8'h3c;
end 13'h19ec:    begin Red = 8'h39;    Green = 8'h1d;    Blue = 8'h43;
end 13'h19ed:    begin Red = 8'h02;    Green = 8'h11;    Blue = 8'h57;
end 13'h19ee:    begin Red = 8'h01;    Green = 8'h01;    Blue = 8'h28;
end 13'h19ef:    begin Red = 8'hfe;    Green = 8'hee;    Blue = 8'hbd;
end 13'h19f0:    begin Red = 8'h7f;    Green = 8'h79;    Blue = 8'h73;
end 13'h19f1:    begin Red = 8'h84;    Green = 8'h7e;    Blue = 8'h78;
end 13'h19f2:    begin Red = 8'h6a;    Green = 8'h8d;    Blue = 8'ha3;
end 13'h19f3:    begin Red = 8'h65;    Green = 8'h89;    Blue = 8'ha0;
end 13'h19f4:    begin Red = 8'h6e;    Green = 8'h65;    Blue = 8'h61;
end 13'h19f5:    begin Red = 8'h3a;    Green = 8'h35;    Blue = 8'h35;
end 13'h19f6:    begin Red = 8'ha0;    Green = 8'haf;    Blue = 8'hb7;
end 13'h19f7:    begin Red = 8'h9e;    Green = 8'hb3;    Blue = 8'hb2;
end 13'h19f8:    begin Red = 8'h90;    Green = 8'h9b;    Blue = 8'ha2;
end 13'h19f9:    begin Red = 8'h9a;    Green = 8'haa;    Blue = 8'hb3;
end 13'h19fa:    begin Red = 8'h7d;    Green = 8'hcc;    Blue = 8'hfd;
end 13'h19fb:    begin Red = 8'h74;    Green = 8'hb9;    Blue = 8'he4;
end 13'h19fc:    begin Red = 8'h4e;    Green = 8'h79;    Blue = 8'hb1;
end 13'h19fd:    begin Red = 8'hf0;    Green = 8'he5;    Blue = 8'he5;
end 13'h19fe:    begin Red = 8'h94;    Green = 8'h92;    Blue = 8'h57;
end 13'h19ff:    begin Red = 8'h79;    Green = 8'h78;    Blue = 8'h42;
end 13'h1a00:    begin Red = 8'h64;    Green = 8'h68;    Blue = 8'h36;
end 13'h1a01:    begin Red = 8'h61;    Green = 8'h60;    Blue = 8'h32;
end 13'h1a02:    begin Red = 8'h50;    Green = 8'h5c;    Blue = 8'h2a;
end 13'h1a03:    begin Red = 8'h63;    Green = 8'h5c;    Blue = 8'h2e;
end 13'h1a04:    begin Red = 8'h42;    Green = 8'h4d;    Blue = 8'h25;
end 13'h1a05:    begin Red = 8'he6;    Green = 8'hd1;    Blue = 8'ha2;
end 13'h1a06:    begin Red = 8'hd7;    Green = 8'hbb;    Blue = 8'h89;
end 13'h1a07:    begin Red = 8'h82;    Green = 8'h8b;    Blue = 8'h9a;
end 13'h1a08:    begin Red = 8'hb2;    Green = 8'hd4;    Blue = 8'hdd;
end 13'h1a09:    begin Red = 8'hb3;    Green = 8'hd9;    Blue = 8'hdc;
end 13'h1a0a:    begin Red = 8'hb8;    Green = 8'hd9;    Blue = 8'hce;
end 13'h1a0b:    begin Red = 8'hb8;    Green = 8'hd6;    Blue = 8'hd4;
end 13'h1a0c:    begin Red = 8'hc5;    Green = 8'h45;    Blue = 8'h42;
end 13'h1a0d:    begin Red = 8'hd3;    Green = 8'hb5;    Blue = 8'h83;
end 13'h1a0e:    begin Red = 8'hef;    Green = 8'hce;    Blue = 8'hab;
end 13'h1a0f:    begin Red = 8'h4c;    Green = 8'h35;    Blue = 8'h2f;
end 13'h1a10:    begin Red = 8'h49;    Green = 8'h34;    Blue = 8'h31;
end 13'h1a11:    begin Red = 8'h4a;    Green = 8'h2e;    Blue = 8'h47;
end 13'h1a12:    begin Red = 8'h51;    Green = 8'h2c;    Blue = 8'h58;
end 13'h1a13:    begin Red = 8'h41;    Green = 8'h24;    Blue = 8'h54;
end 13'h1a14:    begin Red = 8'h3e;    Green = 8'h23;    Blue = 8'h4e;
end 13'h1a15:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'h06;
end 13'h1a16:    begin Red = 8'h4b;    Green = 8'h2a;    Blue = 8'h59;
end 13'h1a17:    begin Red = 8'h47;    Green = 8'h2b;    Blue = 8'h53;
end 13'h1a18:    begin Red = 8'h45;    Green = 8'h29;    Blue = 8'h51;
end 13'h1a19:    begin Red = 8'h42;    Green = 8'h27;    Blue = 8'h52;
end 13'h1a1a:    begin Red = 8'h3d;    Green = 8'h1f;    Blue = 8'h5b;
end 13'h1a1b:    begin Red = 8'h40;    Green = 8'h23;    Blue = 8'h51;
end 13'h1a1c:    begin Red = 8'h3e;    Green = 8'h20;    Blue = 8'h54;
end 13'h1a1d:    begin Red = 8'h7a;    Green = 8'h66;    Blue = 8'h71;
end 13'h1a1e:    begin Red = 8'h72;    Green = 8'h60;    Blue = 8'h6c;
end 13'h1a1f:    begin Red = 8'h01;    Green = 8'he1;    Blue = 8'h5e;
end 13'h1a20:    begin Red = 8'h47;    Green = 8'h2a;    Blue = 8'h58;
end 13'h1a21:    begin Red = 8'h48;    Green = 8'h27;    Blue = 8'h52;
end 13'h1a22:    begin Red = 8'h36;    Green = 8'h1a;    Blue = 8'h4d;
end 13'h1a23:    begin Red = 8'h78;    Green = 8'h65;    Blue = 8'h6b;
end 13'h1a24:    begin Red = 8'h01;    Green = 8'h40;    Blue = 8'h3b;
end 13'h1a25:    begin Red = 8'h50;    Green = 8'h4a;    Blue = 8'h55;
end 13'h1a26:    begin Red = 8'hb3;    Green = 8'ha8;    Blue = 8'h9b;
end 13'h1a27:    begin Red = 8'haf;    Green = 8'ha3;    Blue = 8'h99;
end 13'h1a28:    begin Red = 8'hf1;    Green = 8'he5;    Blue = 8'hce;
end 13'h1a29:    begin Red = 8'h3f;    Green = 8'h3f;    Blue = 8'h3b;
end 13'h1a2a:    begin Red = 8'h59;    Green = 8'h4f;    Blue = 8'h4f;
end 13'h1a2b:    begin Red = 8'h69;    Green = 8'h5e;    Blue = 8'h65;
end 13'h1a2c:    begin Red = 8'hb5;    Green = 8'ha3;    Blue = 8'h83;
end 13'h1a2d:    begin Red = 8'h6a;    Green = 8'h94;    Blue = 8'h42;
end 13'h1a2e:    begin Red = 8'h68;    Green = 8'h92;    Blue = 8'h3e;
end 13'h1a2f:    begin Red = 8'h67;    Green = 8'h90;    Blue = 8'h41;
end 13'h1a30:    begin Red = 8'h69;    Green = 8'h92;    Blue = 8'h46;
end 13'h1a31:    begin Red = 8'h52;    Green = 8'h71;    Blue = 8'h36;
end 13'h1a32:    begin Red = 8'h57;    Green = 8'h70;    Blue = 8'h2f;
end 13'h1a33:    begin Red = 8'h38;    Green = 8'h5d;    Blue = 8'h1a;
end 13'h1a34:    begin Red = 8'hab;    Green = 8'hb0;    Blue = 8'h8d;
end 13'h1a35:    begin Red = 8'h6a;    Green = 8'h62;    Blue = 8'h3b;
end 13'h1a36:    begin Red = 8'h6a;    Green = 8'h71;    Blue = 8'h3e;
end 13'h1a37:    begin Red = 8'h60;    Green = 8'h64;    Blue = 8'h32;
end 13'h1a38:    begin Red = 8'h7f;    Green = 8'h72;    Blue = 8'h4f;
end 13'h1a39:    begin Red = 8'h76;    Green = 8'h6d;    Blue = 8'h44;
end 13'h1a3a:    begin Red = 8'h5f;    Green = 8'h5a;    Blue = 8'h30;
end 13'h1a3b:    begin Red = 8'h48;    Green = 8'h4f;    Blue = 8'h23;
end 13'h1a3c:    begin Red = 8'h49;    Green = 8'h49;    Blue = 8'h25;
end 13'h1a3d:    begin Red = 8'hd9;    Green = 8'hde;    Blue = 8'hbe;
end 13'h1a3e:    begin Red = 8'h99;    Green = 8'h8e;    Blue = 8'h77;
end 13'h1a3f:    begin Red = 8'hd2;    Green = 8'hb4;    Blue = 8'h80;
end 13'h1a40:    begin Red = 8'h8a;    Green = 8'h94;    Blue = 8'h9d;
end 13'h1a41:    begin Red = 8'h04;    Green = 8'h6b;    Blue = 8'h1d;
end 13'h1a42:    begin Red = 8'h10;    Green = 8'h1c;    Blue = 8'h2a;
end 13'h1a43:    begin Red = 8'h1e;    Green = 8'h1c;    Blue = 8'h29;
end 13'h1a44:    begin Red = 8'h1c;    Green = 8'h20;    Blue = 8'h23;
end 13'h1a45:    begin Red = 8'h60;    Green = 8'h75;    Blue = 8'h86;
end 13'h1a46:    begin Red = 8'h08;    Green = 8'h26;    Blue = 8'h14;
end 13'h1a47:    begin Red = 8'he9;    Green = 8'hd3;    Blue = 8'ha4;
end 13'h1a48:    begin Red = 8'hed;    Green = 8'hd0;    Blue = 8'ha4;
end 13'h1a49:    begin Red = 8'h4b;    Green = 8'h2e;    Blue = 8'h40;
end 13'h1a4a:    begin Red = 8'h4f;    Green = 8'h3c;    Blue = 8'h38;
end 13'h1a4b:    begin Red = 8'h51;    Green = 8'h38;    Blue = 8'h3e;
end 13'h1a4c:    begin Red = 8'h54;    Green = 8'h33;    Blue = 8'h4e;
end 13'h1a4d:    begin Red = 8'hc7;    Green = 8'hae;    Blue = 8'h78;
end 13'h1a4e:    begin Red = 8'h54;    Green = 8'h49;    Blue = 8'h33;
end 13'h1a4f:    begin Red = 8'hea;    Green = 8'hf6;    Blue = 8'hd2;
end 13'h1a50:    begin Red = 8'h36;    Green = 8'h26;    Blue = 8'h27;
end 13'h1a51:    begin Red = 8'h02;    Green = 8'h01;    Blue = 8'h2f;
end 13'h1a52:    begin Red = 8'h3b;    Green = 8'h28;    Blue = 8'h24;
end 13'h1a53:    begin Red = 8'h2d;    Green = 8'h24;    Blue = 8'h13;
end 13'h1a54:    begin Red = 8'h23;    Green = 8'h17;    Blue = 8'h17;
end 13'h1a55:    begin Red = 8'h22;    Green = 8'h16;    Blue = 8'h24;
end 13'h1a56:    begin Red = 8'h01;    Green = 8'he1;    Blue = 8'h4b;
end 13'h1a57:    begin Red = 8'h00;    Green = 8'h18;    Blue = 8'hfa;
end 13'h1a58:    begin Red = 8'h27;    Green = 8'h17;    Blue = 8'h22;
end 13'h1a59:    begin Red = 8'h2e;    Green = 8'h23;    Blue = 8'h21;
end 13'h1a5a:    begin Red = 8'h31;    Green = 8'h23;    Blue = 8'h1a;
end 13'h1a5b:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'h04;
end 13'h1a5c:    begin Red = 8'hce;    Green = 8'hb2;    Blue = 8'h80;
end 13'h1a5d:    begin Red = 8'h64;    Green = 8'h5d;    Blue = 8'h5b;
end 13'h1a5e:    begin Red = 8'h5e;    Green = 8'h5f;    Blue = 8'h52;
end 13'h1a5f:    begin Red = 8'h57;    Green = 8'h4f;    Blue = 8'h56;
end 13'h1a60:    begin Red = 8'hb3;    Green = 8'hae;    Blue = 8'ha9;
end 13'h1a61:    begin Red = 8'hba;    Green = 8'hb3;    Blue = 8'had;
end 13'h1a62:    begin Red = 8'hb5;    Green = 8'hb1;    Blue = 8'haf;
end 13'h1a63:    begin Red = 8'ha4;    Green = 8'h9d;    Blue = 8'h98;
end 13'h1a64:    begin Red = 8'hc7;    Green = 8'hc5;    Blue = 8'hbb;
end 13'h1a65:    begin Red = 8'hc1;    Green = 8'hc0;    Blue = 8'hb2;
end 13'h1a66:    begin Red = 8'ha7;    Green = 8'hac;    Blue = 8'ha7;
end 13'h1a67:    begin Red = 8'hc0;    Green = 8'hbd;    Blue = 8'hb4;
end 13'h1a68:    begin Red = 8'hb2;    Green = 8'haa;    Blue = 8'ha9;
end 13'h1a69:    begin Red = 8'h6a;    Green = 8'h8d;    Blue = 8'h4d;
end 13'h1a6a:    begin Red = 8'h00;    Green = 8'h1d;    Blue = 8'h07;
end 13'h1a6b:    begin Red = 8'h02;    Green = 8'haa;    Blue = 8'h17;
end 13'h1a6c:    begin Red = 8'h00;    Green = 8'h07;    Blue = 8'h13;
end 13'h1a6d:    begin Red = 8'h00;    Green = 8'h08;    Blue = 8'h26;
end 13'h1a6e:    begin Red = 8'h49;    Green = 8'h70;    Blue = 8'h2d;
end 13'h1a6f:    begin Red = 8'h3e;    Green = 8'h5e;    Blue = 8'h1d;
end 13'h1a70:    begin Red = 8'hf7;    Green = 8'hea;    Blue = 8'hbd;
end 13'h1a71:    begin Red = 8'hee;    Green = 8'he4;    Blue = 8'hbb;
end 13'h1a72:    begin Red = 8'h06;    Green = 8'h83;    Blue = 8'hda;
end 13'h1a73:    begin Red = 8'h04;    Green = 8'h12;    Blue = 8'h97;
end 13'h1a74:    begin Red = 8'h6f;    Green = 8'h6d;    Blue = 8'h44;
end 13'h1a75:    begin Red = 8'h5c;    Green = 8'h54;    Blue = 8'h2f;
end 13'h1a76:    begin Red = 8'h85;    Green = 8'h92;    Blue = 8'h98;
end 13'h1a77:    begin Red = 8'h63;    Green = 8'h34;    Blue = 8'h48;
end 13'h1a78:    begin Red = 8'h32;    Green = 8'h40;    Blue = 8'h49;
end 13'h1a79:    begin Red = 8'h3b;    Green = 8'h3f;    Blue = 8'h4a;
end 13'h1a7a:    begin Red = 8'h3a;    Green = 8'h39;    Blue = 8'h3f;
end 13'h1a7b:    begin Red = 8'h3e;    Green = 8'h45;    Blue = 8'h4f;
end 13'h1a7c:    begin Red = 8'h7a;    Green = 8'h77;    Blue = 8'h94;
end 13'h1a7d:    begin Red = 8'h69;    Green = 8'h74;    Blue = 8'h7a;
end 13'h1a7e:    begin Red = 8'h7f;    Green = 8'h69;    Blue = 8'h14;
end 13'h1a7f:    begin Red = 8'h4b;    Green = 8'h3a;    Blue = 8'h30;
end 13'h1a80:    begin Red = 8'h4d;    Green = 8'h3a;    Blue = 8'h34;
end 13'h1a81:    begin Red = 8'h4f;    Green = 8'h31;    Blue = 8'h4b;
end 13'h1a82:    begin Red = 8'hea;    Green = 8'hf1;    Blue = 8'hcc;
end 13'h1a83:    begin Red = 8'h34;    Green = 8'h28;    Blue = 8'h36;
end 13'h1a84:    begin Red = 8'h2f;    Green = 8'h26;    Blue = 8'h2b;
end 13'h1a85:    begin Red = 8'h22;    Green = 8'h12;    Blue = 8'h12;
end 13'h1a86:    begin Red = 8'h30;    Green = 8'h23;    Blue = 8'h2a;
end 13'h1a87:    begin Red = 8'h2e;    Green = 8'h20;    Blue = 8'h2f;
end 13'h1a88:    begin Red = 8'h01;    Green = 8'hf1;    Blue = 8'h0b;
end 13'h1a89:    begin Red = 8'h00;    Green = 8'h1c;    Blue = 8'hed;
end 13'h1a8a:    begin Red = 8'h34;    Green = 8'h25;    Blue = 8'h2a;
end 13'h1a8b:    begin Red = 8'h3a;    Green = 8'h29;    Blue = 8'h2f;
end 13'h1a8c:    begin Red = 8'h63;    Green = 8'h5c;    Blue = 8'h60;
end 13'h1a8d:    begin Red = 8'h62;    Green = 8'h5c;    Blue = 8'h66;
end 13'h1a8e:    begin Red = 8'h6d;    Green = 8'h5a;    Blue = 8'h6a;
end 13'h1a8f:    begin Red = 8'h87;    Green = 8'h84;    Blue = 8'h80;
end 13'h1a90:    begin Red = 8'haf;    Green = 8'hac;    Blue = 8'ha5;
end 13'h1a91:    begin Red = 8'hb4;    Green = 8'hab;    Blue = 8'hab;
end 13'h1a92:    begin Red = 8'hb1;    Green = 8'hae;    Blue = 8'ha4;
end 13'h1a93:    begin Red = 8'hac;    Green = 8'ha8;    Blue = 8'ha5;
end 13'h1a94:    begin Red = 8'h6e;    Green = 8'h94;    Blue = 8'h3f;
end 13'h1a95:    begin Red = 8'h02;    Green = 8'hcd;    Blue = 8'h1f;
end 13'h1a96:    begin Red = 8'h01;    Green = 8'h11;    Blue = 8'h2a;
end 13'h1a97:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h2f;
end 13'h1a98:    begin Red = 8'h1c;    Green = 8'h14;    Blue = 8'h11;
end 13'h1a99:    begin Red = 8'h18;    Green = 8'h15;    Blue = 8'h10;
end 13'h1a9a:    begin Red = 8'h01;    Green = 8'h71;    Blue = 8'h4f;
end 13'h1a9b:    begin Red = 8'h01;    Green = 8'h61;    Blue = 8'h3e;
end 13'h1a9c:    begin Red = 8'h01;    Green = 8'hc1;    Blue = 8'h3e;
end 13'h1a9d:    begin Red = 8'h53;    Green = 8'h75;    Blue = 8'h39;
end 13'h1a9e:    begin Red = 8'h44;    Green = 8'h68;    Blue = 8'h28;
end 13'h1a9f:    begin Red = 8'hea;    Green = 8'hdc;    Blue = 8'hb6;
end 13'h1aa0:    begin Red = 8'hed;    Green = 8'hdb;    Blue = 8'hba;
end 13'h1aa1:    begin Red = 8'h7c;    Green = 8'h7b;    Blue = 8'h4b;
end 13'h1aa2:    begin Red = 8'h64;    Green = 8'h6a;    Blue = 8'h3a;
end 13'h1aa3:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'ha4;
end 13'h1aa4:    begin Red = 8'h4d;    Green = 8'h54;    Blue = 8'h2a;
end 13'h1aa5:    begin Red = 8'h85;    Green = 8'h65;    Blue = 8'h18;
end 13'h1aa6:    begin Red = 8'h38;    Green = 8'h41;    Blue = 8'h4a;
end 13'h1aa7:    begin Red = 8'h2d;    Green = 8'h29;    Blue = 8'h37;
end 13'h1aa8:    begin Red = 8'h2b;    Green = 8'h27;    Blue = 8'h35;
end 13'h1aa9:    begin Red = 8'h2d;    Green = 8'h34;    Blue = 8'h3e;
end 13'h1aaa:    begin Red = 8'h69;    Green = 8'h72;    Blue = 8'h81;
end 13'h1aab:    begin Red = 8'h3b;    Green = 8'h3b;    Blue = 8'h47;
end 13'h1aac:    begin Red = 8'h08;    Green = 8'h36;    Blue = 8'h04;
end 13'h1aad:    begin Red = 8'hc3;    Green = 8'hb0;    Blue = 8'h76;
end 13'h1aae:    begin Red = 8'h54;    Green = 8'h40;    Blue = 8'h37;
end 13'h1aaf:    begin Red = 8'h54;    Green = 8'h3c;    Blue = 8'h3c;
end 13'h1ab0:    begin Red = 8'h57;    Green = 8'h37;    Blue = 8'h4c;
end 13'h1ab1:    begin Red = 8'h57;    Green = 8'h36;    Blue = 8'h51;
end 13'h1ab2:    begin Red = 8'hfd;    Green = 8'hf4;    Blue = 8'haf;
end 13'h1ab3:    begin Red = 8'h5b;    Green = 8'h2e;    Blue = 8'h69;
end 13'h1ab4:    begin Red = 8'hce;    Green = 8'hd9;    Blue = 8'hab;
end 13'h1ab5:    begin Red = 8'h49;    Green = 8'h25;    Blue = 8'h62;
end 13'h1ab6:    begin Red = 8'h4b;    Green = 8'h23;    Blue = 8'h5f;
end 13'h1ab7:    begin Red = 8'h01;    Green = 8'he1;    Blue = 8'h3d;
end 13'h1ab8:    begin Red = 8'h00;    Green = 8'h14;    Blue = 8'hf0;
end 13'h1ab9:    begin Red = 8'h55;    Green = 8'h2d;    Blue = 8'h69;
end 13'h1aba:    begin Red = 8'h54;    Green = 8'h2b;    Blue = 8'h67;
end 13'h1abb:    begin Red = 8'h4f;    Green = 8'h27;    Blue = 8'h63;
end 13'h1abc:    begin Red = 8'h47;    Green = 8'h23;    Blue = 8'h60;
end 13'h1abd:    begin Red = 8'h00;    Green = 8'h1b;    Blue = 8'he5;
end 13'h1abe:    begin Red = 8'h4c;    Green = 8'h2a;    Blue = 8'h66;
end 13'h1abf:    begin Red = 8'h51;    Green = 8'h25;    Blue = 8'h60;
end 13'h1ac0:    begin Red = 8'h47;    Green = 8'h24;    Blue = 8'h5a;
end 13'h1ac1:    begin Red = 8'h50;    Green = 8'h23;    Blue = 8'h5e;
end 13'h1ac2:    begin Red = 8'h02;    Green = 8'h60;    Blue = 8'h57;
end 13'h1ac3:    begin Red = 8'h60;    Green = 8'h50;    Blue = 8'h57;
end 13'h1ac4:    begin Red = 8'h68;    Green = 8'h96;    Blue = 8'h68;
end 13'h1ac5:    begin Red = 8'h60;    Green = 8'h51;    Blue = 8'h61;
end 13'h1ac6:    begin Red = 8'h5a;    Green = 8'h52;    Blue = 8'h55;
end 13'h1ac7:    begin Red = 8'h5e;    Green = 8'h3e;    Blue = 8'h25;
end 13'h1ac8:    begin Red = 8'h02;    Green = 8'h87;    Blue = 8'h1a;
end 13'h1ac9:    begin Red = 8'h35;    Green = 8'h24;    Blue = 8'h1d;
end 13'h1aca:    begin Red = 8'h01;    Green = 8'h31;    Blue = 8'h2d;
end 13'h1acb:    begin Red = 8'h01;    Green = 8'h21;    Blue = 8'h1f;
end 13'h1acc:    begin Red = 8'h00;    Green = 8'h0f;    Blue = 8'hec;
end 13'h1acd:    begin Red = 8'h01;    Green = 8'ha1;    Blue = 8'h2f;
end 13'h1ace:    begin Red = 8'h00;    Green = 8'h14;    Blue = 8'hf9;
end 13'h1acf:    begin Red = 8'h01;    Green = 8'hb1;    Blue = 8'h1f;
end 13'h1ad0:    begin Red = 8'h56;    Green = 8'h77;    Blue = 8'h32;
end 13'h1ad1:    begin Red = 8'h5a;    Green = 8'h42;    Blue = 8'h26;
end 13'h1ad2:    begin Red = 8'h8a;    Green = 8'h8a;    Blue = 8'h4e;
end 13'h1ad3:    begin Red = 8'h85;    Green = 8'h82;    Blue = 8'h4f;
end 13'h1ad4:    begin Red = 8'h67;    Green = 8'h6b;    Blue = 8'h39;
end 13'h1ad5:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'hc4;
end 13'h1ad6:    begin Red = 8'h45;    Green = 8'h4c;    Blue = 8'h22;
end 13'h1ad7:    begin Red = 8'he9;    Green = 8'hcd;    Blue = 8'ha8;
end 13'h1ad8:    begin Red = 8'h1e;    Green = 8'h20;    Blue = 8'h2c;
end 13'h1ad9:    begin Red = 8'h95;    Green = 8'ha2;    Blue = 8'haa;
end 13'h1ada:    begin Red = 8'h33;    Green = 8'h2f;    Blue = 8'h3d;
end 13'h1adb:    begin Red = 8'h77;    Green = 8'h7d;    Blue = 8'h8b;
end 13'h1adc:    begin Red = 8'h2b;    Green = 8'h2e;    Blue = 8'h3d;
end 13'h1add:    begin Red = 8'h32;    Green = 8'h34;    Blue = 8'h40;
end 13'h1ade:    begin Red = 8'h07;    Green = 8'hf6;    Blue = 8'h0e;
end 13'h1adf:    begin Red = 8'h08;    Green = 8'h26;    Blue = 8'h06;
end 13'h1ae0:    begin Red = 8'hae;    Green = 8'h98;    Blue = 8'h6f;
end 13'h1ae1:    begin Red = 8'h55;    Green = 8'h3d;    Blue = 8'h39;
end 13'h1ae2:    begin Red = 8'h55;    Green = 8'h39;    Blue = 8'h45;
end 13'h1ae3:    begin Red = 8'hbf;    Green = 8'haa;    Blue = 8'h71;
end 13'h1ae4:    begin Red = 8'hc7;    Green = 8'hd6;    Blue = 8'ha4;
end 13'h1ae5:    begin Red = 8'h4c;    Green = 8'h25;    Blue = 8'h64;
end 13'h1ae6:    begin Red = 8'h00;    Green = 8'h14;    Blue = 8'hd0;
end 13'h1ae7:    begin Red = 8'h51;    Green = 8'h2b;    Blue = 8'h64;
end 13'h1ae8:    begin Red = 8'h38;    Green = 8'h21;    Blue = 8'h71;
end 13'h1ae9:    begin Red = 8'h33;    Green = 8'h22;    Blue = 8'h70;
end 13'h1aea:    begin Red = 8'h2d;    Green = 8'h1c;    Blue = 8'h6a;
end 13'h1aeb:    begin Red = 8'h2f;    Green = 8'h25;    Blue = 8'h6e;
end 13'h1aec:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h58;
end 13'h1aed:    begin Red = 8'h5c;    Green = 8'h58;    Blue = 8'h55;
end 13'h1aee:    begin Red = 8'h62;    Green = 8'ha5;    Blue = 8'h67;
end 13'h1aef:    begin Red = 8'h65;    Green = 8'h51;    Blue = 8'h5c;
end 13'h1af0:    begin Red = 8'hac;    Green = 8'ha9;    Blue = 8'ha0;
end 13'h1af1:    begin Red = 8'h3e;    Green = 8'h35;    Blue = 8'h14;
end 13'h1af2:    begin Red = 8'h3c;    Green = 8'h51;    Blue = 8'h26;
end 13'h1af3:    begin Red = 8'h66;    Green = 8'h93;    Blue = 8'h42;
end 13'h1af4:    begin Red = 8'h00;    Green = 8'h20;    Blue = 8'h0f;
end 13'h1af5:    begin Red = 8'h02;    Green = 8'hac;    Blue = 8'h14;
end 13'h1af6:    begin Red = 8'h00;    Green = 8'h00;    Blue = 8'h04;
end 13'h1af7:    begin Red = 8'h02;    Green = 8'h5b;    Blue = 8'h14;
end 13'h1af8:    begin Red = 8'h00;    Green = 8'h09;    Blue = 8'h56;
end 13'h1af9:    begin Red = 8'h01;    Green = 8'h51;    Blue = 8'h2d;
end 13'h1afa:    begin Red = 8'h17;    Green = 8'h11;    Blue = 8'h13;
end 13'h1afb:    begin Red = 8'h00;    Green = 8'h0a;    Blue = 8'h05;
end 13'h1afc:    begin Red = 8'h45;    Green = 8'h7f;    Blue = 8'h44;
end 13'h1afd:    begin Red = 8'h3f;    Green = 8'h4c;    Blue = 8'h32;
end 13'h1afe:    begin Red = 8'h98;    Green = 8'haf;    Blue = 8'ha7;
end 13'h1aff:    begin Red = 8'h04;    Green = 8'he2;    Blue = 8'hf3;
end 13'h1b00:    begin Red = 8'h8e;    Green = 8'h8b;    Blue = 8'h54;
end 13'h1b01:    begin Red = 8'h06;    Green = 8'h83;    Blue = 8'hcb;
end 13'h1b02:    begin Red = 8'h04;    Green = 8'h42;    Blue = 8'hd4;
end 13'h1b03:    begin Red = 8'h76;    Green = 8'h73;    Blue = 8'h48;
end 13'h1b04:    begin Red = 8'hd2;    Green = 8'hb5;    Blue = 8'h89;
end 13'h1b05:    begin Red = 8'h82;    Green = 8'h67;    Blue = 8'h18;
end 13'h1b06:    begin Red = 8'h81;    Green = 8'h90;    Blue = 8'h97;
end 13'h1b07:    begin Red = 8'h92;    Green = 8'ha7;    Blue = 8'hac;
end 13'h1b08:    begin Red = 8'h40;    Green = 8'h42;    Blue = 8'h4e;
end 13'h1b09:    begin Red = 8'h74;    Green = 8'h77;    Blue = 8'h86;
end 13'h1b0a:    begin Red = 8'h6b;    Green = 8'h6e;    Blue = 8'h7d;
end 13'h1b0b:    begin Red = 8'he7;    Green = 8'hcb;    Blue = 8'ha3;
end 13'h1b0c:    begin Red = 8'h5a;    Green = 8'h42;    Blue = 8'h3e;
end 13'h1b0d:    begin Red = 8'h5c;    Green = 8'h42;    Blue = 8'h43;
end 13'h1b0e:    begin Red = 8'h5d;    Green = 8'h41;    Blue = 8'h40;
end 13'h1b0f:    begin Red = 8'h5c;    Green = 8'h3c;    Blue = 8'h4b;
end 13'h1b10:    begin Red = 8'h5c;    Green = 8'h3a;    Blue = 8'h52;
end 13'h1b11:    begin Red = 8'hfe;    Green = 8'hf0;    Blue = 8'haf;
end 13'h1b12:    begin Red = 8'h5e;    Green = 8'h2d;    Blue = 8'h6f;
end 13'h1b13:    begin Red = 8'h50;    Green = 8'h27;    Blue = 8'h69;
end 13'h1b14:    begin Red = 8'h58;    Green = 8'h2e;    Blue = 8'h6e;
end 13'h1b15:    begin Red = 8'h56;    Green = 8'h2c;    Blue = 8'h6c;
end 13'h1b16:    begin Red = 8'h51;    Green = 8'h2a;    Blue = 8'h6d;
end 13'h1b17:    begin Red = 8'h00;    Green = 8'h19;    Blue = 8'hd1;
end 13'h1b18:    begin Red = 8'h4f;    Green = 8'h2e;    Blue = 8'h67;
end 13'h1b19:    begin Red = 8'hc0;    Green = 8'h3e;    Blue = 8'h31;
end 13'h1b1a:    begin Red = 8'hba;    Green = 8'h41;    Blue = 8'h38;
end 13'h1b1b:    begin Red = 8'hb3;    Green = 8'h3f;    Blue = 8'h32;
end 13'h1b1c:    begin Red = 8'hbf;    Green = 8'h3f;    Blue = 8'h34;
end 13'h1b1d:    begin Red = 8'h49;    Green = 8'h29;    Blue = 8'h6a;
end 13'h1b1e:    begin Red = 8'h02;    Green = 8'hb0;    Blue = 8'h5a;
end 13'h1b1f:    begin Red = 8'hae;    Green = 8'ha8;    Blue = 8'ha2;
end 13'h1b20:    begin Red = 8'h00;    Green = 8'he8;    Blue = 8'h22;
end 13'h1b21:    begin Red = 8'h00;    Green = 8'hdd;    Blue = 8'ha3;
end 13'h1b22:    begin Red = 8'h5d;    Green = 8'h38;    Blue = 8'h32;
end 13'h1b23:    begin Red = 8'h2a;    Green = 8'h19;    Blue = 8'h11;
end 13'h1b24:    begin Red = 8'h2a;    Green = 8'h18;    Blue = 8'h16;
end 13'h1b25:    begin Red = 8'h25;    Green = 8'h15;    Blue = 8'h15;
end 13'h1b26:    begin Red = 8'h50;    Green = 8'h7d;    Blue = 8'h38;
end 13'h1b27:    begin Red = 8'h51;    Green = 8'h75;    Blue = 8'h35;
end 13'h1b28:    begin Red = 8'h39;    Green = 8'h87;    Blue = 8'h49;
end 13'h1b29:    begin Red = 8'h00;    Green = 8'hdf;    Blue = 8'hac;
end 13'h1b2a:    begin Red = 8'h87;    Green = 8'hb2;    Blue = 8'hab;
end 13'h1b2b:    begin Red = 8'hc4;    Green = 8'hb8;    Blue = 8'h9e;
end 13'h1b2c:    begin Red = 8'h04;    Green = 8'hb2;    Blue = 8'hc0;
end 13'h1b2d:    begin Red = 8'h82;    Green = 8'h7a;    Blue = 8'h4b;
end 13'h1b2e:    begin Red = 8'h7d;    Green = 8'h7d;    Blue = 8'h47;
end 13'h1b2f:    begin Red = 8'h55;    Green = 8'h53;    Blue = 8'h20;
end 13'h1b30:    begin Red = 8'h2c;    Green = 8'h3b;    Blue = 8'h3e;
end 13'h1b31:    begin Red = 8'h1a;    Green = 8'h3e;    Blue = 8'h58;
end 13'h1b32:    begin Red = 8'h0b;    Green = 8'hf2;    Blue = 8'h7f;
end 13'h1b33:    begin Red = 8'hb3;    Green = 8'h27;    Blue = 8'h18;
end 13'h1b34:    begin Red = 8'hba;    Green = 8'h2c;    Blue = 8'h16;
end 13'h1b35:    begin Red = 8'hbb;    Green = 8'h2d;    Blue = 8'h19;
end 13'h1b36:    begin Red = 8'hb6;    Green = 8'h28;    Blue = 8'h12;
end 13'h1b37:    begin Red = 8'hba;    Green = 8'h28;    Blue = 8'h19;
end 13'h1b38:    begin Red = 8'hbf;    Green = 8'h28;    Blue = 8'h21;
end 13'h1b39:    begin Red = 8'hc3;    Green = 8'h25;    Blue = 8'h1a;
end 13'h1b3a:    begin Red = 8'hb8;    Green = 8'h25;    Blue = 8'h1b;
end 13'h1b3b:    begin Red = 8'hb9;    Green = 8'h23;    Blue = 8'h22;
end 13'h1b3c:    begin Red = 8'h8d;    Green = 8'h21;    Blue = 8'h15;
end 13'h1b3d:    begin Red = 8'h88;    Green = 8'h19;    Blue = 8'h12;
end 13'h1b3e:    begin Red = 8'h82;    Green = 8'h23;    Blue = 8'h11;
end 13'h1b3f:    begin Red = 8'h5f;    Green = 8'h4c;    Blue = 8'h68;
end 13'h1b40:    begin Red = 8'h56;    Green = 8'h4c;    Blue = 8'h65;
end 13'h1b41:    begin Red = 8'ha5;    Green = 8'h92;    Blue = 8'h68;
end 13'h1b42:    begin Red = 8'h5d;    Green = 8'h47;    Blue = 8'h3c;
end 13'h1b43:    begin Red = 8'h5f;    Green = 8'h3d;    Blue = 8'h55;
end 13'h1b44:    begin Red = 8'hba;    Green = 8'ha5;    Blue = 8'h6e;
end 13'h1b45:    begin Red = 8'h53;    Green = 8'h47;    Blue = 8'h31;
end 13'h1b46:    begin Red = 8'hff;    Green = 8'hee;    Blue = 8'hac;
end 13'h1b47:    begin Red = 8'h46;    Green = 8'h1f;    Blue = 8'h60;
end 13'h1b48:    begin Red = 8'hb7;    Green = 8'hbc;    Blue = 8'h9e;
end 13'h1b49:    begin Red = 8'h38;    Green = 8'h1b;    Blue = 8'h5e;
end 13'h1b4a:    begin Red = 8'h2c;    Green = 8'h1c;    Blue = 8'h5d;
end 13'h1b4b:    begin Red = 8'h35;    Green = 8'h1c;    Blue = 8'h60;
end 13'h1b4c:    begin Red = 8'h3c;    Green = 8'h1f;    Blue = 8'h5f;
end 13'h1b4d:    begin Red = 8'h58;    Green = 8'h2b;    Blue = 8'h70;
end 13'h1b4e:    begin Red = 8'h5b;    Green = 8'h27;    Blue = 8'h6f;
end 13'h1b4f:    begin Red = 8'h2d;    Green = 8'h1e;    Blue = 8'h59;
end 13'h1b50:    begin Red = 8'h36;    Green = 8'h1c;    Blue = 8'h5b;
end 13'h1b51:    begin Red = 8'h32;    Green = 8'h18;    Blue = 8'h57;
end 13'h1b52:    begin Red = 8'h4e;    Green = 8'h29;    Blue = 8'h6c;
end 13'h1b53:    begin Red = 8'h54;    Green = 8'h2d;    Blue = 8'h70;
end 13'h1b54:    begin Red = 8'h1d;    Green = 8'h11;    Blue = 8'h15;
end 13'h1b55:    begin Red = 8'h01;    Green = 8'he1;    Blue = 8'h30;
end 13'h1b56:    begin Red = 8'hb3;    Green = 8'h44;    Blue = 8'h31;
end 13'h1b57:    begin Red = 8'hb8;    Green = 8'h43;    Blue = 8'h39;
end 13'h1b58:    begin Red = 8'hb6;    Green = 8'h42;    Blue = 8'h42;
end 13'h1b59:    begin Red = 8'h58;    Green = 8'h24;    Blue = 8'h77;
end 13'h1b5a:    begin Red = 8'h37;    Green = 8'h17;    Blue = 8'h58;
end 13'h1b5b:    begin Red = 8'h33;    Green = 8'h15;    Blue = 8'h55;
end 13'h1b5c:    begin Red = 8'h3a;    Green = 8'h1d;    Blue = 8'h60;
end 13'h1b5d:    begin Red = 8'h00;    Green = 8'hf2;    Blue = 8'h48;
end 13'h1b5e:    begin Red = 8'h83;    Green = 8'h84;    Blue = 8'h7f;
end 13'h1b5f:    begin Red = 8'h1c;    Green = 8'h5b;    Blue = 8'h87;
end 13'h1b60:    begin Red = 8'h1c;    Green = 8'h5f;    Blue = 8'h96;
end 13'h1b61:    begin Red = 8'h34;    Green = 8'h2c;    Blue = 8'h2a;
end 13'h1b62:    begin Red = 8'h21;    Green = 8'h5d;    Blue = 8'h9b;
end 13'h1b63:    begin Red = 8'h27;    Green = 8'h4f;    Blue = 8'h80;
end 13'h1b64:    begin Red = 8'hb1;    Green = 8'ha1;    Blue = 8'h9b;
end 13'h1b65:    begin Red = 8'haf;    Green = 8'ha2;    Blue = 8'haa;
end 13'h1b66:    begin Red = 8'h00;    Green = 8'hea;    Blue = 8'h03;
end 13'h1b67:    begin Red = 8'h00;    Green = 8'he1;    Blue = 8'h6e;
end 13'h1b68:    begin Red = 8'h68;    Green = 8'h9d;    Blue = 8'h43;
end 13'h1b69:    begin Red = 8'h65;    Green = 8'h46;    Blue = 8'h41;
end 13'h1b6a:    begin Red = 8'h7e;    Green = 8'h5f;    Blue = 8'h4b;
end 13'h1b6b:    begin Red = 8'h74;    Green = 8'h5c;    Blue = 8'h4f;
end 13'h1b6c:    begin Red = 8'h5a;    Green = 8'h51;    Blue = 8'h30;
end 13'h1b6d:    begin Red = 8'h53;    Green = 8'h73;    Blue = 8'h41;
end 13'h1b6e:    begin Red = 8'h4c;    Green = 8'h6a;    Blue = 8'h34;
end 13'h1b6f:    begin Red = 8'h6b;    Green = 8'h91;    Blue = 8'h44;
end 13'h1b70:    begin Red = 8'h4f;    Green = 8'h74;    Blue = 8'h40;
end 13'h1b71:    begin Red = 8'h32;    Green = 8'h8a;    Blue = 8'h4d;
end 13'h1b72:    begin Red = 8'h00;    Green = 8'he4;    Blue = 8'hb6;
end 13'h1b73:    begin Red = 8'h87;    Green = 8'hb0;    Blue = 8'ha2;
end 13'h1b74:    begin Red = 8'hd9;    Green = 8'hcb;    Blue = 8'ha9;
end 13'h1b75:    begin Red = 8'hbd;    Green = 8'hb3;    Blue = 8'h90;
end 13'h1b76:    begin Red = 8'hbd;    Green = 8'hb0;    Blue = 8'h96;
end 13'h1b77:    begin Red = 8'hd7;    Green = 8'haf;    Blue = 8'h74;
end 13'h1b78:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'h61;
end 13'h1b79:    begin Red = 8'h04;    Green = 8'hd2;    Blue = 8'hc0;
end 13'h1b7a:    begin Red = 8'h5c;    Green = 8'h66;    Blue = 8'h34;
end 13'h1b7b:    begin Red = 8'h06;    Green = 8'h53;    Blue = 8'he7;
end 13'h1b7c:    begin Red = 8'hde;    Green = 8'hb8;    Blue = 8'h7a;
end 13'h1b7d:    begin Red = 8'h04;    Green = 8'h62;    Blue = 8'h97;
end 13'h1b7e:    begin Red = 8'h04;    Green = 8'h12;    Blue = 8'hb2;
end 13'h1b7f:    begin Red = 8'h77;    Green = 8'h6f;    Blue = 8'h41;
end 13'h1b80:    begin Red = 8'h62;    Green = 8'h63;    Blue = 8'h39;
end 13'h1b81:    begin Red = 8'h4e;    Green = 8'h49;    Blue = 8'h23;
end 13'h1b82:    begin Red = 8'h05;    Green = 8'h53;    Blue = 8'h67;
end 13'h1b83:    begin Red = 8'hb4;    Green = 8'h94;    Blue = 8'h63;
end 13'h1b84:    begin Red = 8'h86;    Green = 8'h70;    Blue = 8'h58;
end 13'h1b85:    begin Red = 8'h82;    Green = 8'h63;    Blue = 8'h20;
end 13'h1b86:    begin Red = 8'h0c;    Green = 8'h3e;    Blue = 8'h45;
end 13'h1b87:    begin Red = 8'hb9;    Green = 8'h22;    Blue = 8'h19;
end 13'h1b88:    begin Red = 8'hba;    Green = 8'h2b;    Blue = 8'h1d;
end 13'h1b89:    begin Red = 8'hbd;    Green = 8'h27;    Blue = 8'h16;
end 13'h1b8a:    begin Red = 8'hbf;    Green = 8'h27;    Blue = 8'h1a;
end 13'h1b8b:    begin Red = 8'h83;    Green = 8'h21;    Blue = 8'h18;
end 13'h1b8c:    begin Red = 8'h8a;    Green = 8'h1d;    Blue = 8'h16;
end 13'h1b8d:    begin Red = 8'h89;    Green = 8'h23;    Blue = 8'h14;
end 13'h1b8e:    begin Red = 8'h58;    Green = 8'h50;    Blue = 8'h68;
end 13'h1b8f:    begin Red = 8'h5f;    Green = 8'h4a;    Blue = 8'h6b;
end 13'h1b90:    begin Red = 8'hcb;    Green = 8'hbd;    Blue = 8'h8e;
end 13'h1b91:    begin Red = 8'h5b;    Green = 8'h50;    Blue = 8'h3e;
end 13'h1b92:    begin Red = 8'h5f;    Green = 8'h48;    Blue = 8'h40;
end 13'h1b93:    begin Red = 8'h5f;    Green = 8'h45;    Blue = 8'h44;
end 13'h1b94:    begin Red = 8'h5e;    Green = 8'h44;    Blue = 8'h47;
end 13'h1b95:    begin Red = 8'h60;    Green = 8'h3f;    Blue = 8'h50;
end 13'h1b96:    begin Red = 8'hc9;    Green = 8'haf;    Blue = 8'h7c;
end 13'h1b97:    begin Red = 8'hec;    Green = 8'hf7;    Blue = 8'hc8;
end 13'h1b98:    begin Red = 8'h36;    Green = 8'h17;    Blue = 8'h50;
end 13'h1b99:    begin Red = 8'h34;    Green = 8'h1a;    Blue = 8'h63;
end 13'h1b9a:    begin Red = 8'h33;    Green = 8'h1d;    Blue = 8'h5d;
end 13'h1b9b:    begin Red = 8'h01;    Green = 8'h81;    Blue = 8'h10;
end 13'h1b9c:    begin Red = 8'h42;    Green = 8'h24;    Blue = 8'h58;
end 13'h1b9d:    begin Red = 8'h3a;    Green = 8'h1c;    Blue = 8'h5c;
end 13'h1b9e:    begin Red = 8'h2e;    Green = 8'h19;    Blue = 8'h54;
end 13'h1b9f:    begin Red = 8'h4f;    Green = 8'h2f;    Blue = 8'h6e;
end 13'h1ba0:    begin Red = 8'h58;    Green = 8'h24;    Blue = 8'h62;
end 13'h1ba1:    begin Red = 8'h1b;    Green = 8'h17;    Blue = 8'h18;
end 13'h1ba2:    begin Red = 8'hc0;    Green = 8'h3f;    Blue = 8'h3a;
end 13'h1ba3:    begin Red = 8'hb8;    Green = 8'h3f;    Blue = 8'h2c;
end 13'h1ba4:    begin Red = 8'h58;    Green = 8'h2d;    Blue = 8'h63;
end 13'h1ba5:    begin Red = 8'h35;    Green = 8'h1b;    Blue = 8'h58;
end 13'h1ba6:    begin Red = 8'h31;    Green = 8'h17;    Blue = 8'h54;
end 13'h1ba7:    begin Red = 8'hff;    Green = 8'he2;    Blue = 8'hb6;
end 13'h1ba8:    begin Red = 8'h60;    Green = 8'h5b;    Blue = 8'h5e;
end 13'h1ba9:    begin Red = 8'h87;    Green = 8'h7f;    Blue = 8'h7d;
end 13'h1baa:    begin Red = 8'h20;    Green = 8'h53;    Blue = 8'h82;
end 13'h1bab:    begin Red = 8'h2b;    Green = 8'h54;    Blue = 8'h82;
end 13'h1bac:    begin Red = 8'h00;    Green = 8'hf3;    Blue = 8'h03;
end 13'h1bad:    begin Red = 8'h00;    Green = 8'he4;    Blue = 8'h4c;
end 13'h1bae:    begin Red = 8'h6a;    Green = 8'h92;    Blue = 8'h4c;
end 13'h1baf:    begin Red = 8'h70;    Green = 8'ha2;    Blue = 8'h5d;
end 13'h1bb0:    begin Red = 8'h6f;    Green = 8'h5b;    Blue = 8'h52;
end 13'h1bb1:    begin Red = 8'h70;    Green = 8'h5e;    Blue = 8'h46;
end 13'h1bb2:    begin Red = 8'h72;    Green = 8'h5a;    Blue = 8'h50;
end 13'h1bb3:    begin Red = 8'h6d;    Green = 8'h58;    Blue = 8'h47;
end 13'h1bb4:    begin Red = 8'h58;    Green = 8'h4e;    Blue = 8'h33;
end 13'h1bb5:    begin Red = 8'h6c;    Green = 8'h96;    Blue = 8'h44;
end 13'h1bb6:    begin Red = 8'h2f;    Green = 8'h89;    Blue = 8'h43;
end 13'h1bb7:    begin Red = 8'h0d;    Green = 8'ha8;    Blue = 8'h13;
end 13'h1bb8:    begin Red = 8'h8e;    Green = 8'hb6;    Blue = 8'hae;
end 13'h1bb9:    begin Red = 8'hd7;    Green = 8'hca;    Blue = 8'ha7;
end 13'h1bba:    begin Red = 8'hf1;    Green = 8'hc3;    Blue = 8'h85;
end 13'h1bbb:    begin Red = 8'h02;    Green = 8'he1;    Blue = 8'h45;
end 13'h1bbc:    begin Red = 8'h59;    Green = 8'h62;    Blue = 8'h33;
end 13'h1bbd:    begin Red = 8'h54;    Green = 8'h5d;    Blue = 8'h30;
end 13'h1bbe:    begin Red = 8'h06;    Green = 8'hb4;    Blue = 8'h2c;
end 13'h1bbf:    begin Red = 8'he1;    Green = 8'hbf;    Blue = 8'h7f;
end 13'h1bc0:    begin Red = 8'h04;    Green = 8'h52;    Blue = 8'h73;
end 13'h1bc1:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'ha2;
end 13'h1bc2:    begin Red = 8'h7a;    Green = 8'h6d;    Blue = 8'h41;
end 13'h1bc3:    begin Red = 8'h66;    Green = 8'h67;    Blue = 8'h3d;
end 13'h1bc4:    begin Red = 8'h51;    Green = 8'h4c;    Blue = 8'h24;
end 13'h1bc5:    begin Red = 8'h41;    Green = 8'h4a;    Blue = 8'h1f;
end 13'h1bc6:    begin Red = 8'h8b;    Green = 8'h6b;    Blue = 8'h42;
end 13'h1bc7:    begin Red = 8'hcb;    Green = 8'hae;    Blue = 8'h84;
end 13'h1bc8:    begin Red = 8'he6;    Green = 8'hc8;    Blue = 8'ha4;
end 13'h1bc9:    begin Red = 8'hd6;    Green = 8'hab;    Blue = 8'h89;
end 13'h1bca:    begin Red = 8'h74;    Green = 8'h82;    Blue = 8'h61;
end 13'h1bcb:    begin Red = 8'h52;    Green = 8'h55;    Blue = 8'h76;
end 13'h1bcc:    begin Red = 8'h4e;    Green = 8'h4f;    Blue = 8'h7b;
end 13'h1bcd:    begin Red = 8'h4b;    Green = 8'h4e;    Blue = 8'h77;
end 13'h1bce:    begin Red = 8'h56;    Green = 8'h55;    Blue = 8'h74;
end 13'h1bcf:    begin Red = 8'h54;    Green = 8'h52;    Blue = 8'h79;
end 13'h1bd0:    begin Red = 8'h28;    Green = 8'h29;    Blue = 8'h3b;
end 13'h1bd1:    begin Red = 8'h33;    Green = 8'h31;    Blue = 8'h49;
end 13'h1bd2:    begin Red = 8'h16;    Green = 8'h33;    Blue = 8'h53;
end 13'h1bd3:    begin Red = 8'hb2;    Green = 8'h2a;    Blue = 8'h10;
end 13'h1bd4:    begin Red = 8'h8e;    Green = 8'h1b;    Blue = 8'h14;
end 13'h1bd5:    begin Red = 8'h87;    Green = 8'h20;    Blue = 8'h19;
end 13'h1bd6:    begin Red = 8'h60;    Green = 8'h51;    Blue = 8'h66;
end 13'h1bd7:    begin Red = 8'h5c;    Green = 8'h4e;    Blue = 8'h67;
end 13'h1bd8:    begin Red = 8'hcf;    Green = 8'had;    Blue = 8'h87;
end 13'h1bd9:    begin Red = 8'h62;    Green = 8'h4b;    Blue = 8'h3b;
end 13'h1bda:    begin Red = 8'h61;    Green = 8'h48;    Blue = 8'h44;
end 13'h1bdb:    begin Red = 8'h62;    Green = 8'h44;    Blue = 8'h46;
end 13'h1bdc:    begin Red = 8'h63;    Green = 8'h42;    Blue = 8'h53;
end 13'h1bdd:    begin Red = 8'h62;    Green = 8'h41;    Blue = 8'h56;
end 13'h1bde:    begin Red = 8'hb4;    Green = 8'ha1;    Blue = 8'h67;
end 13'h1bdf:    begin Red = 8'ha0;    Green = 8'h93;    Blue = 8'h69;
end 13'h1be0:    begin Red = 8'hc9;    Green = 8'hb1;    Blue = 8'h83;
end 13'h1be1:    begin Red = 8'hde;    Green = 8'hc9;    Blue = 8'h9e;
end 13'h1be2:    begin Red = 8'hee;    Green = 8'hf7;    Blue = 8'hd5;
end 13'h1be3:    begin Red = 8'hb4;    Green = 8'h43;    Blue = 8'h35;
end 13'h1be4:    begin Red = 8'hbb;    Green = 8'h3f;    Blue = 8'h33;
end 13'h1be5:    begin Red = 8'h4e;    Green = 8'h47;    Blue = 8'h34;
end 13'h1be6:    begin Red = 8'h15;    Green = 8'h4e;    Blue = 8'h93;
end 13'h1be7:    begin Red = 8'h21;    Green = 8'h16;    Blue = 8'h1c;
end 13'h1be8:    begin Red = 8'h1d;    Green = 8'h19;    Blue = 8'h1a;
end 13'h1be9:    begin Red = 8'h02;    Green = 8'h21;    Blue = 8'h8c;
end 13'h1bea:    begin Red = 8'h24;    Green = 8'h1a;    Blue = 8'h11;
end 13'h1beb:    begin Red = 8'h1c;    Green = 8'h1c;    Blue = 8'h14;
end 13'h1bec:    begin Red = 8'h22;    Green = 8'h1a;    Blue = 8'h18;
end 13'h1bed:    begin Red = 8'h1e;    Green = 8'h1d;    Blue = 8'h18;
end 13'h1bee:    begin Red = 8'h02;    Green = 8'h41;    Blue = 8'h7e;
end 13'h1bef:    begin Red = 8'h07;    Green = 8'h49;    Blue = 8'h86;
end 13'h1bf0:    begin Red = 8'h3e;    Green = 8'h5a;    Blue = 8'h20;
end 13'h1bf1:    begin Red = 8'h4c;    Green = 8'h64;    Blue = 8'h34;
end 13'h1bf2:    begin Red = 8'h7b;    Green = 8'had;    Blue = 8'h56;
end 13'h1bf3:    begin Red = 8'h52;    Green = 8'hbc;    Blue = 8'hf0;
end 13'h1bf4:    begin Red = 8'h00;    Green = 8'h1b;    Blue = 8'h99;
end 13'h1bf5:    begin Red = 8'h78;    Green = 8'h69;    Blue = 8'h6c;
end 13'h1bf6:    begin Red = 8'had;    Green = 8'ha3;    Blue = 8'h84;
end 13'h1bf7:    begin Red = 8'hae;    Green = 8'ha5;    Blue = 8'h81;
end 13'h1bf8:    begin Red = 8'hbb;    Green = 8'haf;    Blue = 8'h92;
end 13'h1bf9:    begin Red = 8'hcf;    Green = 8'haf;    Blue = 8'h7c;
end 13'h1bfa:    begin Red = 8'h03;    Green = 8'h21;    Blue = 8'h04;
end 13'h1bfb:    begin Red = 8'h04;    Green = 8'hd2;    Blue = 8'hb0;
end 13'h1bfc:    begin Red = 8'h06;    Green = 8'hd3;    Blue = 8'h9a;
end 13'h1bfd:    begin Red = 8'hf3;    Green = 8'hda;    Blue = 8'ha1;
end 13'h1bfe:    begin Red = 8'hdb;    Green = 8'hbb;    Blue = 8'h80;
end 13'h1bff:    begin Red = 8'hdc;    Green = 8'hb7;    Blue = 8'h82;
end 13'h1c00:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'h70;
end 13'h1c01:    begin Red = 8'h42;    Green = 8'h3d;    Blue = 8'h17;
end 13'h1c02:    begin Red = 8'h3f;    Green = 8'h46;    Blue = 8'h24;
end 13'h1c03:    begin Red = 8'h3b;    Green = 8'h42;    Blue = 8'h20;
end 13'h1c04:    begin Red = 8'h3e;    Green = 8'h43;    Blue = 8'h1b;
end 13'h1c05:    begin Red = 8'h05;    Green = 8'h33;    Blue = 8'h34;
end 13'h1c06:    begin Red = 8'he2;    Green = 8'hd0;    Blue = 8'ha0;
end 13'h1c07:    begin Red = 8'hd2;    Green = 8'hce;    Blue = 8'ha1;
end 13'h1c08:    begin Red = 8'hec;    Green = 8'hef;    Blue = 8'hc2;
end 13'h1c09:    begin Red = 8'h6a;    Green = 8'h8b;    Blue = 8'h5c;
end 13'h1c0a:    begin Red = 8'h0d;    Green = 8'h01;    Blue = 8'h5c;
end 13'h1c0b:    begin Red = 8'h57;    Green = 8'h4c;    Blue = 8'h77;
end 13'h1c0c:    begin Red = 8'h44;    Green = 8'h4b;    Blue = 8'h79;
end 13'h1c0d:    begin Red = 8'h50;    Green = 8'h50;    Blue = 8'h68;
end 13'h1c0e:    begin Red = 8'h53;    Green = 8'h51;    Blue = 8'h76;
end 13'h1c0f:    begin Red = 8'h5c;    Green = 8'h5b;    Blue = 8'h7d;
end 13'h1c10:    begin Red = 8'hb1;    Green = 8'h24;    Blue = 8'h12;
end 13'h1c11:    begin Red = 8'hb3;    Green = 8'h2e;    Blue = 8'h1d;
end 13'h1c12:    begin Red = 8'h08;    Green = 8'h31;    Blue = 8'h99;
end 13'h1c13:    begin Red = 8'h76;    Green = 8'h1e;    Blue = 8'h1c;
end 13'h1c14:    begin Red = 8'h5d;    Green = 8'h58;    Blue = 8'h78;
end 13'h1c15:    begin Red = 8'h58;    Green = 8'h51;    Blue = 8'h7d;
end 13'h1c16:    begin Red = 8'he0;    Green = 8'hc3;    Blue = 8'h99;
end 13'h1c17:    begin Red = 8'h3b;    Green = 8'h31;    Blue = 8'h25;
end 13'h1c18:    begin Red = 8'ha8;    Green = 8'h91;    Blue = 8'h65;
end 13'h1c19:    begin Red = 8'hbd;    Green = 8'ha6;    Blue = 8'h74;
end 13'h1c1a:    begin Red = 8'h62;    Green = 8'h55;    Blue = 8'h21;
end 13'h1c1b:    begin Red = 8'h67;    Green = 8'h55;    Blue = 8'h27;
end 13'h1c1c:    begin Red = 8'h5f;    Green = 8'h49;    Blue = 8'h3b;
end 13'h1c1d:    begin Red = 8'h62;    Green = 8'h44;    Blue = 8'h4c;
end 13'h1c1e:    begin Red = 8'hfb;    Green = 8'he8;    Blue = 8'hc0;
end 13'h1c1f:    begin Red = 8'h00;    Green = 8'h07;    Blue = 8'h32;
end 13'h1c20:    begin Red = 8'h00;    Green = 8'h0c;    Blue = 8'h10;
end 13'h1c21:    begin Red = 8'h00;    Green = 8'h0c;    Blue = 8'h21;
end 13'h1c22:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'h45;
end 13'h1c23:    begin Red = 8'hbc;    Green = 8'h26;    Blue = 8'h27;
end 13'h1c24:    begin Red = 8'hc4;    Green = 8'h31;    Blue = 8'h27;
end 13'h1c25:    begin Red = 8'hd4;    Green = 8'h3f;    Blue = 8'h38;
end 13'h1c26:    begin Red = 8'hba;    Green = 8'h2a;    Blue = 8'h22;
end 13'h1c27:    begin Red = 8'haa;    Green = 8'h2b;    Blue = 8'h22;
end 13'h1c28:    begin Red = 8'h00;    Green = 8'h08;    Blue = 8'h41;
end 13'h1c29:    begin Red = 8'h65;    Green = 8'h59;    Blue = 8'h5a;
end 13'h1c2a:    begin Red = 8'h04;    Green = 8'h48;    Blue = 8'h89;
end 13'h1c2b:    begin Red = 8'h26;    Green = 8'h54;    Blue = 8'h92;
end 13'h1c2c:    begin Red = 8'h00;    Green = 8'h1f;    Blue = 8'hc0;
end 13'h1c2d:    begin Red = 8'h00;    Green = 8'h24;    Blue = 8'ha0;
end 13'h1c2e:    begin Red = 8'h00;    Green = 8'h25;    Blue = 8'hb0;
end 13'h1c2f:    begin Red = 8'h00;    Green = 8'h1f;    Blue = 8'h61;
end 13'h1c30:    begin Red = 8'h00;    Green = 8'h27;    Blue = 8'h90;
end 13'h1c31:    begin Red = 8'h00;    Green = 8'h16;    Blue = 8'h30;
end 13'h1c32:    begin Red = 8'h00;    Green = 8'h23;    Blue = 8'h73;
end 13'h1c33:    begin Red = 8'h00;    Green = 8'h20;    Blue = 8'h01;
end 13'h1c34:    begin Red = 8'h00;    Green = 8'h29;    Blue = 8'h00;
end 13'h1c35:    begin Red = 8'h00;    Green = 8'h22;    Blue = 8'h30;
end 13'h1c36:    begin Red = 8'h1d;    Green = 8'h56;    Blue = 8'h8b;
end 13'h1c37:    begin Red = 8'h77;    Green = 8'h75;    Blue = 8'h68;
end 13'h1c38:    begin Red = 8'hb3;    Green = 8'ha3;    Blue = 8'ha8;
end 13'h1c39:    begin Red = 8'h42;    Green = 8'h59;    Blue = 8'h21;
end 13'h1c3a:    begin Red = 8'h54;    Green = 8'h73;    Blue = 8'h37;
end 13'h1c3b:    begin Red = 8'h4e;    Green = 8'h69;    Blue = 8'h32;
end 13'h1c3c:    begin Red = 8'h4b;    Green = 8'h67;    Blue = 8'h36;
end 13'h1c3d:    begin Red = 8'h78;    Green = 8'h6c;    Blue = 8'h78;
end 13'h1c3e:    begin Red = 8'h90;    Green = 8'h85;    Blue = 8'h91;
end 13'h1c3f:    begin Red = 8'h8e;    Green = 8'h8a;    Blue = 8'h7a;
end 13'h1c40:    begin Red = 8'h90;    Green = 8'h85;    Blue = 8'h8c;
end 13'h1c41:    begin Red = 8'he2;    Green = 8'hc2;    Blue = 8'h8f;
end 13'h1c42:    begin Red = 8'hef;    Green = 8'hd3;    Blue = 8'ha1;
end 13'h1c43:    begin Red = 8'heb;    Green = 8'hc8;    Blue = 8'h8e;
end 13'h1c44:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'h25;
end 13'h1c45:    begin Red = 8'h04;    Green = 8'h82;    Blue = 8'hc0;
end 13'h1c46:    begin Red = 8'h70;    Green = 8'h6e;    Blue = 8'h3b;
end 13'h1c47:    begin Red = 8'h58;    Green = 8'h55;    Blue = 8'h28;
end 13'h1c48:    begin Red = 8'h48;    Green = 8'h4e;    Blue = 8'h2a;
end 13'h1c49:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'h98;
end 13'h1c4a:    begin Red = 8'hf8;    Green = 8'hd9;    Blue = 8'ha0;
end 13'h1c4b:    begin Red = 8'hc2;    Green = 8'ha4;    Blue = 8'h6e;
end 13'h1c4c:    begin Red = 8'h03;    Green = 8'hc2;    Blue = 8'h91;
end 13'h1c4d:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h83;
end 13'h1c4e:    begin Red = 8'h3d;    Green = 8'h44;    Blue = 8'h25;
end 13'h1c4f:    begin Red = 8'h3b;    Green = 8'h3f;    Blue = 8'h1e;
end 13'h1c50:    begin Red = 8'h05;    Green = 8'h73;    Blue = 8'h78;
end 13'h1c51:    begin Red = 8'hc1;    Green = 8'ha5;    Blue = 8'h76;
end 13'h1c52:    begin Red = 8'hc2;    Green = 8'ha5;    Blue = 8'h7b;
end 13'h1c53:    begin Red = 8'he0;    Green = 8'hca;    Blue = 8'h9b;
end 13'h1c54:    begin Red = 8'he3;    Green = 8'he9;    Blue = 8'hbd;
end 13'h1c55:    begin Red = 8'hb8;    Green = 8'h2c;    Blue = 8'h13;
end 13'h1c56:    begin Red = 8'h0d;    Green = 8'h01;    Blue = 8'hc3;
end 13'h1c57:    begin Red = 8'h51;    Green = 8'h54;    Blue = 8'h73;
end 13'h1c58:    begin Red = 8'h4f;    Green = 8'h54;    Blue = 8'h7a;
end 13'h1c59:    begin Red = 8'h31;    Green = 8'h32;    Blue = 8'h44;
end 13'h1c5a:    begin Red = 8'h32;    Green = 8'h32;    Blue = 8'h4e;
end 13'h1c5b:    begin Red = 8'h83;    Green = 8'h1a;    Blue = 8'h17;
end 13'h1c5c:    begin Red = 8'h83;    Green = 8'h1c;    Blue = 8'h13;
end 13'h1c5d:    begin Red = 8'h87;    Green = 8'h20;    Blue = 8'h11;
end 13'h1c5e:    begin Red = 8'hf4;    Green = 8'he9;    Blue = 8'hbc;
end 13'h1c5f:    begin Red = 8'hdb;    Green = 8'hbf;    Blue = 8'h97;
end 13'h1c60:    begin Red = 8'hb9;    Green = 8'ha2;    Blue = 8'h6c;
end 13'h1c61:    begin Red = 8'h40;    Green = 8'h2b;    Blue = 8'h63;
end 13'h1c62:    begin Red = 8'h3d;    Green = 8'h28;    Blue = 8'h61;
end 13'h1c63:    begin Red = 8'h62;    Green = 8'h4b;    Blue = 8'h43;
end 13'h1c64:    begin Red = 8'h61;    Green = 8'h47;    Blue = 8'h4a;
end 13'h1c65:    begin Red = 8'h60;    Green = 8'h46;    Blue = 8'h51;
end 13'h1c66:    begin Red = 8'hb0;    Green = 8'h9f;    Blue = 8'h67;
end 13'h1c67:    begin Red = 8'h9d;    Green = 8'h8f;    Blue = 8'h68;
end 13'h1c68:    begin Red = 8'hc1;    Green = 8'ha8;    Blue = 8'h80;
end 13'h1c69:    begin Red = 8'hda;    Green = 8'hb5;    Blue = 8'h8b;
end 13'h1c6a:    begin Red = 8'hc5;    Green = 8'ha5;    Blue = 8'h7e;
end 13'h1c6b:    begin Red = 8'h3f;    Green = 8'h6b;    Blue = 8'h9b;
end 13'h1c6c:    begin Red = 8'h36;    Green = 8'h43;    Blue = 8'h73;
end 13'h1c6d:    begin Red = 8'hff;    Green = 8'hfd;    Blue = 8'hf8;
end 13'h1c6e:    begin Red = 8'h00;    Green = 8'h31;    Blue = 8'h6f;
end 13'h1c6f:    begin Red = 8'h25;    Green = 8'h56;    Blue = 8'h90;
end 13'h1c70:    begin Red = 8'h26;    Green = 8'h56;    Blue = 8'h86;
end 13'h1c71:    begin Red = 8'h21;    Green = 8'h52;    Blue = 8'h7b;
end 13'h1c72:    begin Red = 8'h1e;    Green = 8'h6e;    Blue = 8'hb3;
end 13'h1c73:    begin Red = 8'h25;    Green = 8'h6a;    Blue = 8'hb5;
end 13'h1c74:    begin Red = 8'h25;    Green = 8'h6a;    Blue = 8'had;
end 13'h1c75:    begin Red = 8'h28;    Green = 8'hfd;    Blue = 8'hff;
end 13'h1c76:    begin Red = 8'h2a;    Green = 8'hfa;    Blue = 8'hfc;
end 13'h1c77:    begin Red = 8'h25;    Green = 8'hf6;    Blue = 8'hfa;
end 13'h1c78:    begin Red = 8'h22;    Green = 8'hf8;    Blue = 8'hf8;
end 13'h1c79:    begin Red = 8'h24;    Green = 8'h2f;    Blue = 8'h71;
end 13'h1c7a:    begin Red = 8'h23;    Green = 8'h57;    Blue = 8'h89;
end 13'h1c7b:    begin Red = 8'h25;    Green = 8'h58;    Blue = 8'h8d;
end 13'h1c7c:    begin Red = 8'h43;    Green = 8'h66;    Blue = 8'h8a;
end 13'h1c7d:    begin Red = 8'h67;    Green = 8'h93;    Blue = 8'h48;
end 13'h1c7e:    begin Red = 8'h3e;    Green = 8'h5a;    Blue = 8'h31;
end 13'h1c7f:    begin Red = 8'h56;    Green = 8'h77;    Blue = 8'h40;
end 13'h1c80:    begin Red = 8'h59;    Green = 8'h72;    Blue = 8'h39;
end 13'h1c81:    begin Red = 8'h87;    Green = 8'h85;    Blue = 8'h86;
end 13'h1c82:    begin Red = 8'hd8;    Green = 8'hc9;    Blue = 8'haf;
end 13'h1c83:    begin Red = 8'h02;    Green = 8'hc1;    Blue = 8'h30;
end 13'h1c84:    begin Red = 8'h04;    Green = 8'h73;    Blue = 8'h00;
end 13'h1c85:    begin Red = 8'h06;    Green = 8'h44;    Blue = 8'h1b;
end 13'h1c86:    begin Red = 8'h4f;    Green = 8'h48;    Blue = 8'h2b;
end 13'h1c87:    begin Red = 8'h71;    Green = 8'h69;    Blue = 8'h3b;
end 13'h1c88:    begin Red = 8'h4b;    Green = 8'h46;    Blue = 8'h1e;
end 13'h1c89:    begin Red = 8'h05;    Green = 8'h43;    Blue = 8'h36;
end 13'h1c8a:    begin Red = 8'hbb;    Green = 8'h25;    Blue = 8'h17;
end 13'h1c8b:    begin Red = 8'hbd;    Green = 8'h29;    Blue = 8'h1d;
end 13'h1c8c:    begin Red = 8'hb5;    Green = 8'h2d;    Blue = 8'h17;
end 13'h1c8d:    begin Red = 8'h8f;    Green = 8'h23;    Blue = 8'h16;
end 13'h1c8e:    begin Red = 8'h09;    Green = 8'hb2;    Blue = 8'h1a;
end 13'h1c8f:    begin Red = 8'h94;    Green = 8'h20;    Blue = 8'h13;
end 13'h1c90:    begin Red = 8'ha0;    Green = 8'h20;    Blue = 8'h13;
end 13'h1c91:    begin Red = 8'h96;    Green = 8'h1f;    Blue = 8'h1b;
end 13'h1c92:    begin Red = 8'h99;    Green = 8'h20;    Blue = 8'h18;
end 13'h1c93:    begin Red = 8'h99;    Green = 8'h1f;    Blue = 8'h12;
end 13'h1c94:    begin Red = 8'hb2;    Green = 8'h29;    Blue = 8'h16;
end 13'h1c95:    begin Red = 8'hbf;    Green = 8'h21;    Blue = 8'h18;
end 13'h1c96:    begin Red = 8'hb7;    Green = 8'h29;    Blue = 8'h1f;
end 13'h1c97:    begin Red = 8'hc4;    Green = 8'h28;    Blue = 8'h1c;
end 13'h1c98:    begin Red = 8'h84;    Green = 8'h1d;    Blue = 8'h16;
end 13'h1c99:    begin Red = 8'hff;    Green = 8'h91;    Blue = 8'h1d;
end 13'h1c9a:    begin Red = 8'hfb;    Green = 8'h79;    Blue = 8'h25;
end 13'h1c9b:    begin Red = 8'hfe;    Green = 8'h81;    Blue = 8'h24;
end 13'h1c9c:    begin Red = 8'hf6;    Green = 8'h7e;    Blue = 8'h1f;
end 13'h1c9d:    begin Red = 8'hff;    Green = 8'h7f;    Blue = 8'h22;
end 13'h1c9e:    begin Red = 8'hc9;    Green = 8'ha4;    Blue = 8'h70;
end 13'h1c9f:    begin Red = 8'h56;    Green = 8'h48;    Blue = 8'h3b;
end 13'h1ca0:    begin Red = 8'hb2;    Green = 8'ha6;    Blue = 8'h74;
end 13'h1ca1:    begin Red = 8'h5d;    Green = 8'h52;    Blue = 8'h32;
end 13'h1ca2:    begin Red = 8'h5f;    Green = 8'h4d;    Blue = 8'h39;
end 13'h1ca3:    begin Red = 8'h63;    Green = 8'h4b;    Blue = 8'h3f;
end 13'h1ca4:    begin Red = 8'haa;    Green = 8'h9e;    Blue = 8'h6c;
end 13'h1ca5:    begin Red = 8'hd9;    Green = 8'hc2;    Blue = 8'h96;
end 13'h1ca6:    begin Red = 8'hc3;    Green = 8'haa;    Blue = 8'h82;
end 13'h1ca7:    begin Red = 8'hc0;    Green = 8'hca;    Blue = 8'hac;
end 13'h1ca8:    begin Red = 8'hbe;    Green = 8'ha6;    Blue = 8'h82;
end 13'h1ca9:    begin Red = 8'h5c;    Green = 8'h5c;    Blue = 8'h62;
end 13'h1caa:    begin Red = 8'h6a;    Green = 8'h51;    Blue = 8'h50;
end 13'h1cab:    begin Red = 8'h23;    Green = 8'h6e;    Blue = 8'hb1;
end 13'h1cac:    begin Red = 8'h1f;    Green = 8'h6a;    Blue = 8'had;
end 13'h1cad:    begin Red = 8'h28;    Green = 8'h6b;    Blue = 8'hb9;
end 13'h1cae:    begin Red = 8'h1c;    Green = 8'h6e;    Blue = 8'haa;
end 13'h1caf:    begin Red = 8'h25;    Green = 8'h65;    Blue = 8'hbc;
end 13'h1cb0:    begin Red = 8'h30;    Green = 8'hf7;    Blue = 8'hfe;
end 13'h1cb1:    begin Red = 8'h1f;    Green = 8'hfd;    Blue = 8'hff;
end 13'h1cb2:    begin Red = 8'h24;    Green = 8'h5d;    Blue = 8'h8a;
end 13'h1cb3:    begin Red = 8'hf7;    Green = 8'hff;    Blue = 8'hff;
end 13'h1cb4:    begin Red = 8'hfa;    Green = 8'hf9;    Blue = 8'hfe;
end 13'h1cb5:    begin Red = 8'h23;    Green = 8'hf6;    Blue = 8'hf0;
end 13'h1cb6:    begin Red = 8'h82;    Green = 8'h84;    Blue = 8'h78;
end 13'h1cb7:    begin Red = 8'h80;    Green = 8'h7e;    Blue = 8'h7a;
end 13'h1cb8:    begin Red = 8'h45;    Green = 8'h5a;    Blue = 8'h31;
end 13'h1cb9:    begin Red = 8'h47;    Green = 8'h62;    Blue = 8'h2f;
end 13'h1cba:    begin Red = 8'h72;    Green = 8'h94;    Blue = 8'h48;
end 13'h1cbb:    begin Red = 8'h6f;    Green = 8'h92;    Blue = 8'h52;
end 13'h1cbc:    begin Red = 8'h75;    Green = 8'h5c;    Blue = 8'h3d;
end 13'h1cbd:    begin Red = 8'h71;    Green = 8'h5c;    Blue = 8'h3f;
end 13'h1cbe:    begin Red = 8'h62;    Green = 8'h45;    Blue = 8'h33;
end 13'h1cbf:    begin Red = 8'h51;    Green = 8'h72;    Blue = 8'h3d;
end 13'h1cc0:    begin Red = 8'h57;    Green = 8'h75;    Blue = 8'h43;
end 13'h1cc1:    begin Red = 8'h4c;    Green = 8'h66;    Blue = 8'h39;
end 13'h1cc2:    begin Red = 8'h5f;    Green = 8'h76;    Blue = 8'h40;
end 13'h1cc3:    begin Red = 8'hd5;    Green = 8'hcb;    Blue = 8'haa;
end 13'h1cc4:    begin Red = 8'hdb;    Green = 8'hd0;    Blue = 8'hab;
end 13'h1cc5:    begin Red = 8'h04;    Green = 8'h93;    Blue = 8'h15;
end 13'h1cc6:    begin Red = 8'h56;    Green = 8'h4d;    Blue = 8'h2e;
end 13'h1cc7:    begin Red = 8'h76;    Green = 8'h7a;    Blue = 8'h3f;
end 13'h1cc8:    begin Red = 8'h63;    Green = 8'h6b;    Blue = 8'h32;
end 13'h1cc9:    begin Red = 8'h5c;    Green = 8'h64;    Blue = 8'h2b;
end 13'h1cca:    begin Red = 8'h54;    Green = 8'h5b;    Blue = 8'h27;
end 13'h1ccb:    begin Red = 8'h6d;    Green = 8'h6b;    Blue = 8'h38;
end 13'h1ccc:    begin Red = 8'h58;    Green = 8'h5a;    Blue = 8'h32;
end 13'h1ccd:    begin Red = 8'h4f;    Green = 8'h43;    Blue = 8'h1d;
end 13'h1cce:    begin Red = 8'h3f;    Green = 8'h4e;    Blue = 8'h23;
end 13'h1ccf:    begin Red = 8'h64;    Green = 8'h92;    Blue = 8'h6b;
end 13'h1cd0:    begin Red = 8'hb6;    Green = 8'h24;    Blue = 8'h17;
end 13'h1cd1:    begin Red = 8'hbe;    Green = 8'h2c;    Blue = 8'h1f;
end 13'h1cd2:    begin Red = 8'hce;    Green = 8'h28;    Blue = 8'h1a;
end 13'h1cd3:    begin Red = 8'hd4;    Green = 8'h28;    Blue = 8'h14;
end 13'h1cd4:    begin Red = 8'h0c;    Green = 8'h21;    Blue = 8'h30;
end 13'h1cd5:    begin Red = 8'h0c;    Green = 8'hf6;    Blue = 8'h10;
end 13'h1cd6:    begin Red = 8'h00;    Green = 8'hd5;    Blue = 8'h20;
end 13'h1cd7:    begin Red = 8'h9c;    Green = 8'h20;    Blue = 8'h16;
end 13'h1cd8:    begin Red = 8'h96;    Green = 8'h26;    Blue = 8'h10;
end 13'h1cd9:    begin Red = 8'ha0;    Green = 8'h1c;    Blue = 8'h1a;
end 13'h1cda:    begin Red = 8'h08;    Green = 8'he1;    Blue = 8'he8;
end 13'h1cdb:    begin Red = 8'h09;    Green = 8'h12;    Blue = 8'h1d;
end 13'h1cdc:    begin Red = 8'hb1;    Green = 8'h2e;    Blue = 8'h1a;
end 13'h1cdd:    begin Red = 8'h0b;    Green = 8'hb2;    Blue = 8'hab;
end 13'h1cde:    begin Red = 8'hcd;    Green = 8'h24;    Blue = 8'h11;
end 13'h1cdf:    begin Red = 8'hda;    Green = 8'h28;    Blue = 8'h1a;
end 13'h1ce0:    begin Red = 8'h0b;    Green = 8'he1;    Blue = 8'h10;
end 13'h1ce1:    begin Red = 8'h00;    Green = 8'hc6;    Blue = 8'hf0;
end 13'h1ce2:    begin Red = 8'h00;    Green = 8'hd4;    Blue = 8'h00;
end 13'h1ce3:    begin Red = 8'hb6;    Green = 8'h26;    Blue = 8'h1d;
end 13'h1ce4:    begin Red = 8'h7a;    Green = 8'h1b;    Blue = 8'h19;
end 13'h1ce5:    begin Red = 8'hfb;    Green = 8'ha5;    Blue = 8'h2e;
end 13'h1ce6:    begin Red = 8'hff;    Green = 8'h95;    Blue = 8'h1c;
end 13'h1ce7:    begin Red = 8'hf8;    Green = 8'h80;    Blue = 8'h21;
end 13'h1ce8:    begin Red = 8'hbb;    Green = 8'hbb;    Blue = 8'h95;
end 13'h1ce9:    begin Red = 8'hc3;    Green = 8'ha2;    Blue = 8'h81;
end 13'h1cea:    begin Red = 8'h45;    Green = 8'h23;    Blue = 8'h3b;
end 13'h1ceb:    begin Red = 8'h4c;    Green = 8'h4c;    Blue = 8'h54;
end 13'h1cec:    begin Red = 8'h64;    Green = 8'h44;    Blue = 8'h4f;
end 13'h1ced:    begin Red = 8'h4f;    Green = 8'h43;    Blue = 8'h33;
end 13'h1cee:    begin Red = 8'hbc;    Green = 8'ha3;    Blue = 8'h7b;
end 13'h1cef:    begin Red = 8'h48;    Green = 8'h43;    Blue = 8'h30;
end 13'h1cf0:    begin Red = 8'he0;    Green = 8'hc3;    Blue = 8'ha1;
end 13'h1cf1:    begin Red = 8'h61;    Green = 8'h56;    Blue = 8'h61;
end 13'h1cf2:    begin Red = 8'h21;    Green = 8'h5a;    Blue = 8'h87;
end 13'h1cf3:    begin Red = 8'h21;    Green = 8'h6c;    Blue = 8'hbd;
end 13'h1cf4:    begin Red = 8'h23;    Green = 8'h70;    Blue = 8'hc2;
end 13'h1cf5:    begin Red = 8'h22;    Green = 8'h6e;    Blue = 8'hb9;
end 13'h1cf6:    begin Red = 8'h24;    Green = 8'h65;    Blue = 8'hb5;
end 13'h1cf7:    begin Red = 8'h1c;    Green = 8'h6c;    Blue = 8'hb5;
end 13'h1cf8:    begin Red = 8'h22;    Green = 8'h60;    Blue = 8'hb5;
end 13'h1cf9:    begin Red = 8'h1b;    Green = 8'h4a;    Blue = 8'ha2;
end 13'h1cfa:    begin Red = 8'h1d;    Green = 8'hfc;    Blue = 8'hf9;
end 13'h1cfb:    begin Red = 8'hfb;    Green = 8'hfe;    Blue = 8'hff;
end 13'h1cfc:    begin Red = 8'h1f;    Green = 8'hf1;    Blue = 8'he4;
end 13'h1cfd:    begin Red = 8'h7d;    Green = 8'h79;    Blue = 8'h77;
end 13'h1cfe:    begin Red = 8'h81;    Green = 8'h7b;    Blue = 8'h79;
end 13'h1cff:    begin Red = 8'h4a;    Green = 8'h5f;    Blue = 8'h34;
end 13'h1d00:    begin Red = 8'h46;    Green = 8'h6f;    Blue = 8'h37;
end 13'h1d01:    begin Red = 8'h74;    Green = 8'ha0;    Blue = 8'h51;
end 13'h1d02:    begin Red = 8'h75;    Green = 8'ha5;    Blue = 8'h51;
end 13'h1d03:    begin Red = 8'h6f;    Green = 8'hae;    Blue = 8'h53;
end 13'h1d04:    begin Red = 8'h5c;    Green = 8'h43;    Blue = 8'h3c;
end 13'h1d05:    begin Red = 8'h70;    Green = 8'h5f;    Blue = 8'h4b;
end 13'h1d06:    begin Red = 8'h7a;    Green = 8'h5e;    Blue = 8'h48;
end 13'h1d07:    begin Red = 8'h60;    Green = 8'h40;    Blue = 8'h33;
end 13'h1d08:    begin Red = 8'h5c;    Green = 8'h85;    Blue = 8'h4b;
end 13'h1d09:    begin Red = 8'h4e;    Green = 8'h75;    Blue = 8'h32;
end 13'h1d0a:    begin Red = 8'h55;    Green = 8'h80;    Blue = 8'h38;
end 13'h1d0b:    begin Red = 8'h55;    Green = 8'h83;    Blue = 8'h43;
end 13'h1d0c:    begin Red = 8'hd3;    Green = 8'hc5;    Blue = 8'ha0;
end 13'h1d0d:    begin Red = 8'hd2;    Green = 8'hc6;    Blue = 8'ha5;
end 13'h1d0e:    begin Red = 8'h05;    Green = 8'h02;    Blue = 8'h84;
end 13'h1d0f:    begin Red = 8'h63;    Green = 8'h6c;    Blue = 8'h3f;
end 13'h1d10:    begin Red = 8'h61;    Green = 8'h6b;    Blue = 8'h39;
end 13'h1d11:    begin Red = 8'h52;    Green = 8'h62;    Blue = 8'h31;
end 13'h1d12:    begin Red = 8'h4e;    Green = 8'h61;    Blue = 8'h34;
end 13'h1d13:    begin Red = 8'h06;    Green = 8'hb3;    Blue = 8'ha2;
end 13'h1d14:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h53;
end 13'h1d15:    begin Red = 8'h40;    Green = 8'h58;    Blue = 8'h26;
end 13'h1d16:    begin Red = 8'h3c;    Green = 8'h56;    Blue = 8'h27;
end 13'h1d17:    begin Red = 8'h41;    Green = 8'h4f;    Blue = 8'h2b;
end 13'h1d18:    begin Red = 8'h3e;    Green = 8'h50;    Blue = 8'h2a;
end 13'h1d19:    begin Red = 8'h05;    Green = 8'h73;    Blue = 8'h1d;
end 13'h1d1a:    begin Red = 8'hb8;    Green = 8'h25;    Blue = 8'h13;
end 13'h1d1b:    begin Red = 8'hbf;    Green = 8'h2c;    Blue = 8'h18;
end 13'h1d1c:    begin Red = 8'h0f;    Green = 8'h15;    Blue = 8'h13;
end 13'h1d1d:    begin Red = 8'h90;    Green = 8'h8f;    Blue = 8'h7b;
end 13'h1d1e:    begin Red = 8'h25;    Green = 8'hee;    Blue = 8'hf8;
end 13'h1d1f:    begin Red = 8'h40;    Green = 8'hdd;    Blue = 8'hff;
end 13'h1d20:    begin Red = 8'h9b;    Green = 8'h23;    Blue = 8'h15;
end 13'h1d21:    begin Red = 8'h9c;    Green = 8'h21;    Blue = 8'h11;
end 13'h1d22:    begin Red = 8'hbb;    Green = 8'h24;    Blue = 8'h1d;
end 13'h1d23:    begin Red = 8'h00;    Green = 8'ha1;    Blue = 8'h5f;
end 13'h1d24:    begin Red = 8'h26;    Green = 8'h14;    Blue = 8'h10;
end 13'h1d25:    begin Red = 8'h9d;    Green = 8'h78;    Blue = 8'h66;
end 13'h1d26:    begin Red = 8'h3d;    Green = 8'he0;    Blue = 8'hff;
end 13'h1d27:    begin Red = 8'h07;    Green = 8'hb1;    Blue = 8'hef;
end 13'h1d28:    begin Red = 8'hf8;    Green = 8'h7d;    Blue = 8'h1d;
end 13'h1d29:    begin Red = 8'hd5;    Green = 8'hbb;    Blue = 8'h96;
end 13'h1d2a:    begin Red = 8'h58;    Green = 8'h4b;    Blue = 8'h29;
end 13'h1d2b:    begin Red = 8'hbe;    Green = 8'ha1;    Blue = 8'h75;
end 13'h1d2c:    begin Red = 8'h23;    Green = 8'h54;    Blue = 8'h8c;
end 13'h1d2d:    begin Red = 8'h28;    Green = 8'h59;    Blue = 8'h84;
end 13'h1d2e:    begin Red = 8'h1d;    Green = 8'h54;    Blue = 8'ha4;
end 13'h1d2f:    begin Red = 8'h30;    Green = 8'hf2;    Blue = 8'hfb;
end 13'h1d30:    begin Red = 8'h1f;    Green = 8'h56;    Blue = 8'h7d;
end 13'h1d31:    begin Red = 8'h21;    Green = 8'h6b;    Blue = 8'hb2;
end 13'h1d32:    begin Red = 8'h26;    Green = 8'hf8;    Blue = 8'hf5;
end 13'h1d33:    begin Red = 8'h24;    Green = 8'hfc;    Blue = 8'hf1;
end 13'h1d34:    begin Red = 8'h23;    Green = 8'hfe;    Blue = 8'hfa;
end 13'h1d35:    begin Red = 8'ha5;    Green = 8'ha0;    Blue = 8'h99;
end 13'h1d36:    begin Red = 8'h40;    Green = 8'h28;    Blue = 8'h1c;
end 13'h1d37:    begin Red = 8'h47;    Green = 8'h3c;    Blue = 8'h20;
end 13'h1d38:    begin Red = 8'h48;    Green = 8'h3d;    Blue = 8'h1d;
end 13'h1d39:    begin Red = 8'h46;    Green = 8'h28;    Blue = 8'h1d;
end 13'h1d3a:    begin Red = 8'h6e;    Green = 8'h93;    Blue = 8'h46;
end 13'h1d3b:    begin Red = 8'h2e;    Green = 8'h1b;    Blue = 8'h21;
end 13'h1d3c:    begin Red = 8'h28;    Green = 8'h15;    Blue = 8'h1b;
end 13'h1d3d:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'h9f;
end 13'h1d3e:    begin Red = 8'h4f;    Green = 8'h81;    Blue = 8'h38;
end 13'h1d3f:    begin Red = 8'h51;    Green = 8'h6f;    Blue = 8'h31;
end 13'h1d40:    begin Red = 8'h46;    Green = 8'h3a;    Blue = 8'h22;
end 13'h1d41:    begin Red = 8'h4a;    Green = 8'h3f;    Blue = 8'h1f;
end 13'h1d42:    begin Red = 8'h5d;    Green = 8'h85;    Blue = 8'h46;
end 13'h1d43:    begin Red = 8'h55;    Green = 8'h74;    Blue = 8'h31;
end 13'h1d44:    begin Red = 8'h80;    Green = 8'h78;    Blue = 8'h7b;
end 13'h1d45:    begin Red = 8'h02;    Green = 8'hd1;    Blue = 8'h40;
end 13'h1d46:    begin Red = 8'h04;    Green = 8'hc2;    Blue = 8'hc5;
end 13'h1d47:    begin Red = 8'h07;    Green = 8'h24;    Blue = 8'h49;
end 13'h1d48:    begin Red = 8'h06;    Green = 8'h83;    Blue = 8'he4;
end 13'h1d49:    begin Red = 8'h06;    Green = 8'h73;    Blue = 8'he6;
end 13'h1d4a:    begin Red = 8'h06;    Green = 8'hd3;    Blue = 8'hfd;
end 13'h1d4b:    begin Red = 8'hea;    Green = 8'hbb;    Blue = 8'h85;
end 13'h1d4c:    begin Red = 8'hbd;    Green = 8'h94;    Blue = 8'h5c;
end 13'h1d4d:    begin Red = 8'h06;    Green = 8'h43;    Blue = 8'hc8;
end 13'h1d4e:    begin Red = 8'h04;    Green = 8'hb1;    Blue = 8'h90;
end 13'h1d4f:    begin Red = 8'h05;    Green = 8'h93;    Blue = 8'h36;
end 13'h1d50:    begin Red = 8'h00;    Green = 8'h13;    Blue = 8'h17;
end 13'h1d51:    begin Red = 8'h08;    Green = 8'h81;    Blue = 8'h8d;
end 13'h1d52:    begin Red = 8'h7a;    Green = 8'h1c;    Blue = 8'h10;
end 13'h1d53:    begin Red = 8'h14;    Green = 8'h14;    Blue = 8'h14;
end 13'h1d54:    begin Red = 8'h29;    Green = 8'h16;    Blue = 8'h12;
end 13'h1d55:    begin Red = 8'h00;    Green = 8'h10;    Blue = 8'h30;
end 13'h1d56:    begin Red = 8'ha4;    Green = 8'h7a;    Blue = 8'h64;
end 13'h1d57:    begin Red = 8'h7c;    Green = 8'h23;    Blue = 8'h11;
end 13'h1d58:    begin Red = 8'h79;    Green = 8'h20;    Blue = 8'h12;
end 13'h1d59:    begin Red = 8'h7b;    Green = 8'h1d;    Blue = 8'h13;
end 13'h1d5a:    begin Red = 8'h09;    Green = 8'h41;    Blue = 8'haf;
end 13'h1d5b:    begin Red = 8'h05;    Green = 8'h15;    Blue = 8'h15;
end 13'h1d5c:    begin Red = 8'h34;    Green = 8'h2b;    Blue = 8'h22;
end 13'h1d5d:    begin Red = 8'h48;    Green = 8'h1d;    Blue = 8'h38;
end 13'h1d5e:    begin Red = 8'h00;    Green = 8'hc5;    Blue = 8'h15;
end 13'h1d5f:    begin Red = 8'h01;    Green = 8'h03;    Blue = 8'h1f;
end 13'h1d60:    begin Red = 8'h98;    Green = 8'h86;    Blue = 8'h60;
end 13'h1d61:    begin Red = 8'h63;    Green = 8'h57;    Blue = 8'h3f;
end 13'h1d62:    begin Red = 8'h4f;    Green = 8'h3f;    Blue = 8'h32;
end 13'h1d63:    begin Red = 8'hb5;    Green = 8'h9c;    Blue = 8'h74;
end 13'h1d64:    begin Red = 8'hcf;    Green = 8'hb9;    Blue = 8'h92;
end 13'h1d65:    begin Red = 8'h24;    Green = 8'h5a;    Blue = 8'h80;
end 13'h1d66:    begin Red = 8'h00;    Green = 8'h0d;    Blue = 8'h0a;
end 13'h1d67:    begin Red = 8'h27;    Green = 8'h50;    Blue = 8'h8e;
end 13'h1d68:    begin Red = 8'h22;    Green = 8'h51;    Blue = 8'h7f;
end 13'h1d69:    begin Red = 8'h1d;    Green = 8'h52;    Blue = 8'h7c;
end 13'h1d6a:    begin Red = 8'h1d;    Green = 8'h30;    Blue = 8'h6b;
end 13'h1d6b:    begin Red = 8'h26;    Green = 8'h27;    Blue = 8'h68;
end 13'h1d6c:    begin Red = 8'ha2;    Green = 8'h9c;    Blue = 8'h94;
end 13'h1d6d:    begin Red = 8'h4f;    Green = 8'h3b;    Blue = 8'h16;
end 13'h1d6e:    begin Red = 8'h44;    Green = 8'h2a;    Blue = 8'h13;
end 13'h1d6f:    begin Red = 8'h3e;    Green = 8'h31;    Blue = 8'h1e;
end 13'h1d70:    begin Red = 8'h4d;    Green = 8'h41;    Blue = 8'h27;
end 13'h1d71:    begin Red = 8'h4b;    Green = 8'h42;    Blue = 8'h1b;
end 13'h1d72:    begin Red = 8'h47;    Green = 8'h2c;    Blue = 8'h19;
end 13'h1d73:    begin Red = 8'h47;    Green = 8'h3b;    Blue = 8'h25;
end 13'h1d74:    begin Red = 8'h37;    Green = 8'h30;    Blue = 8'h1d;
end 13'h1d75:    begin Red = 8'h00;    Green = 8'h0f;    Blue = 8'h6b;
end 13'h1d76:    begin Red = 8'h00;    Green = 8'h16;    Blue = 8'h03;
end 13'h1d77:    begin Red = 8'h00;    Green = 8'h0e;    Blue = 8'ha0;
end 13'h1d78:    begin Red = 8'h00;    Green = 8'h06;    Blue = 8'h0b;
end 13'h1d79:    begin Red = 8'hcb;    Green = 8'hbf;    Blue = 8'ha0;
end 13'h1d7a:    begin Red = 8'hc5;    Green = 8'hb9;    Blue = 8'h98;
end 13'h1d7b:    begin Red = 8'hc4;    Green = 8'h99;    Blue = 8'h62;
end 13'h1d7c:    begin Red = 8'h00;    Green = 8'h11;    Blue = 8'h20;
end 13'h1d7d:    begin Red = 8'h02;    Green = 8'h71;    Blue = 8'h70;
end 13'h1d7e:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'h23;
end 13'h1d7f:    begin Red = 8'h03;    Green = 8'ha2;    Blue = 8'h12;
end 13'h1d80:    begin Red = 8'h03;    Green = 8'ha1;    Blue = 8'hf1;
end 13'h1d81:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h01;
end 13'h1d82:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h10;
end 13'h1d83:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h23;
end 13'h1d84:    begin Red = 8'h02;    Green = 8'h41;    Blue = 8'h52;
end 13'h1d85:    begin Red = 8'h03;    Green = 8'h62;    Blue = 8'h40;
end 13'h1d86:    begin Red = 8'h03;    Green = 8'h02;    Blue = 8'h00;
end 13'h1d87:    begin Red = 8'h03;    Green = 8'h31;    Blue = 8'h90;
end 13'h1d88:    begin Red = 8'h03;    Green = 8'h61;    Blue = 8'hd0;
end 13'h1d89:    begin Red = 8'h02;    Green = 8'hf1;    Blue = 8'ha0;
end 13'h1d8a:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'h90;
end 13'h1d8b:    begin Red = 8'hbd;    Green = 8'h94;    Blue = 8'h66;
end 13'h1d8c:    begin Red = 8'ha5;    Green = 8'h9c;    Blue = 8'h83;
end 13'h1d8d:    begin Red = 8'h13;    Green = 8'h18;    Blue = 8'h14;
end 13'h1d8e:    begin Red = 8'h88;    Green = 8'h1c;    Blue = 8'h10;
end 13'h1d8f:    begin Red = 8'h86;    Green = 8'h1e;    Blue = 8'h13;
end 13'h1d90:    begin Red = 8'h14;    Green = 8'h15;    Blue = 8'h1a;
end 13'h1d91:    begin Red = 8'h02;    Green = 8'hd1;    Blue = 8'hbd;
end 13'h1d92:    begin Red = 8'h2d;    Green = 8'h1a;    Blue = 8'h14;
end 13'h1d93:    begin Red = 8'ha3;    Green = 8'ha8;    Blue = 8'h94;
end 13'h1d94:    begin Red = 8'h99;    Green = 8'h26;    Blue = 8'h14;
end 13'h1d95:    begin Red = 8'h81;    Green = 8'h21;    Blue = 8'h13;
end 13'h1d96:    begin Red = 8'h9b;    Green = 8'h1c;    Blue = 8'h15;
end 13'h1d97:    begin Red = 8'h31;    Green = 8'h15;    Blue = 8'h12;
end 13'h1d98:    begin Red = 8'h02;    Green = 8'ha1;    Blue = 8'h6f;
end 13'h1d99:    begin Red = 8'hfe;    Green = 8'hdb;    Blue = 8'hb3;
end 13'h1d9a:    begin Red = 8'hb7;    Green = 8'h9f;    Blue = 8'h71;
end 13'h1d9b:    begin Red = 8'hb4;    Green = 8'ha4;    Blue = 8'h71;
end 13'h1d9c:    begin Red = 8'h46;    Green = 8'h27;    Blue = 8'h37;
end 13'h1d9d:    begin Red = 8'h19;    Green = 8'h11;    Blue = 8'h1e;
end 13'h1d9e:    begin Red = 8'h01;    Green = 8'hbf;    Blue = 8'h1d;
end 13'h1d9f:    begin Red = 8'h5c;    Green = 8'h45;    Blue = 8'h3f;
end 13'h1da0:    begin Red = 8'hdb;    Green = 8'he4;    Blue = 8'hc4;
end 13'h1da1:    begin Red = 8'hba;    Green = 8'h9b;    Blue = 8'h6f;
end 13'h1da2:    begin Red = 8'hd1;    Green = 8'hbd;    Blue = 8'h8b;
end 13'h1da3:    begin Red = 8'h24;    Green = 8'h53;    Blue = 8'h89;
end 13'h1da4:    begin Red = 8'h27;    Green = 8'h57;    Blue = 8'h7f;
end 13'h1da5:    begin Red = 8'h10;    Green = 8'h12;    Blue = 8'h27;
end 13'h1da6:    begin Red = 8'h10;    Green = 8'h14;    Blue = 8'h2f;
end 13'h1da7:    begin Red = 8'h01;    Green = 8'h6d;    Blue = 8'h2a;
end 13'h1da8:    begin Red = 8'h21;    Green = 8'h53;    Blue = 8'h90;
end 13'h1da9:    begin Red = 8'h1c;    Green = 8'h53;    Blue = 8'h89;
end 13'h1daa:    begin Red = 8'h22;    Green = 8'h56;    Blue = 8'h85;
end 13'h1dab:    begin Red = 8'h22;    Green = 8'h19;    Blue = 8'h14;
end 13'h1dac:    begin Red = 8'h55;    Green = 8'h40;    Blue = 8'h21;
end 13'h1dad:    begin Red = 8'h3d;    Green = 8'h2e;    Blue = 8'h31;
end 13'h1dae:    begin Red = 8'h41;    Green = 8'h31;    Blue = 8'h34;
end 13'h1daf:    begin Red = 8'h49;    Green = 8'h3c;    Blue = 8'h19;
end 13'h1db0:    begin Red = 8'h4c;    Green = 8'h36;    Blue = 8'h21;
end 13'h1db1:    begin Red = 8'h3d;    Green = 8'h2f;    Blue = 8'h22;
end 13'h1db2:    begin Red = 8'h36;    Green = 8'h2e;    Blue = 8'h17;
end 13'h1db3:    begin Red = 8'h20;    Green = 8'h19;    Blue = 8'h11;
end 13'h1db4:    begin Red = 8'hc3;    Green = 8'hb7;    Blue = 8'h9b;
end 13'h1db5:    begin Red = 8'hc8;    Green = 8'h9c;    Blue = 8'h5b;
end 13'h1db6:    begin Red = 8'h02;    Green = 8'hf1;    Blue = 8'hb3;
end 13'h1db7:    begin Red = 8'h04;    Green = 8'h72;    Blue = 8'h40;
end 13'h1db8:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'h60;
end 13'h1db9:    begin Red = 8'h03;    Green = 8'he2;    Blue = 8'h77;
end 13'h1dba:    begin Red = 8'hf3;    Green = 8'hc1;    Blue = 8'h84;
end 13'h1dbb:    begin Red = 8'hd3;    Green = 8'h9f;    Blue = 8'h66;
end 13'h1dbc:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'h50;
end 13'h1dbd:    begin Red = 8'h02;    Green = 8'h91;    Blue = 8'h84;
end 13'h1dbe:    begin Red = 8'h03;    Green = 8'hd2;    Blue = 8'h70;
end 13'h1dbf:    begin Red = 8'h03;    Green = 8'h92;    Blue = 8'h70;
end 13'h1dc0:    begin Red = 8'h03;    Green = 8'hc2;    Blue = 8'h13;
end 13'h1dc1:    begin Red = 8'h00;    Green = 8'h15;    Blue = 8'h12;
end 13'h1dc2:    begin Red = 8'h03;    Green = 8'hb2;    Blue = 8'h24;
end 13'h1dc3:    begin Red = 8'h03;    Green = 8'h61;    Blue = 8'hf0;
end 13'h1dc4:    begin Red = 8'h03;    Green = 8'h71;    Blue = 8'he0;
end 13'h1dc5:    begin Red = 8'h03;    Green = 8'h22;    Blue = 8'h21;
end 13'h1dc6:    begin Red = 8'hc7;    Green = 8'h94;    Blue = 8'h65;
end 13'h1dc7:    begin Red = 8'h43;    Green = 8'hb3;    Blue = 8'hfb;
end 13'h1dc8:    begin Red = 8'h43;    Green = 8'h9a;    Blue = 8'hea;
end 13'h1dc9:    begin Red = 8'h00;    Green = 8'h25;    Blue = 8'h01;
end 13'h1dca:    begin Red = 8'h2e;    Green = 8'h15;    Blue = 8'h10;
end 13'h1dcb:    begin Red = 8'h00;    Green = 8'h2d;    Blue = 8'h01;
end 13'h1dcc:    begin Red = 8'h38;    Green = 8'h97;    Blue = 8'heb;
end 13'h1dcd:    begin Red = 8'h32;    Green = 8'h12;    Blue = 8'h15;
end 13'h1dce:    begin Red = 8'h02;    Green = 8'h31;    Blue = 8'h36;
end 13'h1dcf:    begin Red = 8'h02;    Green = 8'hc1;    Blue = 8'h55;
end 13'h1dd0:    begin Red = 8'hd4;    Green = 8'hd0;    Blue = 8'ha3;
end 13'h1dd1:    begin Red = 8'hdb;    Green = 8'hca;    Blue = 8'h9f;
end 13'h1dd2:    begin Red = 8'hd5;    Green = 8'hcc;    Blue = 8'ha5;
end 13'h1dd3:    begin Red = 8'hd4;    Green = 8'hcd;    Blue = 8'h9f;
end 13'h1dd4:    begin Red = 8'h53;    Green = 8'h48;    Blue = 8'h36;
end 13'h1dd5:    begin Red = 8'h20;    Green = 8'h10;    Blue = 8'h1d;
end 13'h1dd6:    begin Red = 8'h01;    Green = 8'hbd;    Blue = 8'h24;
end 13'h1dd7:    begin Red = 8'h02;    Green = 8'h0f;    Blue = 8'h1f;
end 13'h1dd8:    begin Red = 8'h1e;    Green = 8'h10;    Blue = 8'h21;
end 13'h1dd9:    begin Red = 8'h49;    Green = 8'h3c;    Blue = 8'h36;
end 13'h1dda:    begin Red = 8'he2;    Green = 8'hd6;    Blue = 8'hac;
end 13'h1ddb:    begin Red = 8'he5;    Green = 8'hda;    Blue = 8'ha2;
end 13'h1ddc:    begin Red = 8'hcd;    Green = 8'hc0;    Blue = 8'h89;
end 13'h1ddd:    begin Red = 8'hc6;    Green = 8'hc3;    Blue = 8'h90;
end 13'h1dde:    begin Red = 8'hcb;    Green = 8'hc0;    Blue = 8'h93;
end 13'h1ddf:    begin Red = 8'h42;    Green = 8'h2a;    Blue = 8'h26;
end 13'h1de0:    begin Red = 8'h3d;    Green = 8'h30;    Blue = 8'h27;
end 13'h1de1:    begin Red = 8'h3e;    Green = 8'h2b;    Blue = 8'h24;
end 13'h1de2:    begin Red = 8'h01;    Green = 8'h5e;    Blue = 8'h1e;
end 13'h1de3:    begin Red = 8'h14;    Green = 8'h11;    Blue = 8'h2c;
end 13'h1de4:    begin Red = 8'h1a;    Green = 8'h19;    Blue = 8'h38;
end 13'h1de5:    begin Red = 8'h1c;    Green = 8'h16;    Blue = 8'h38;
end 13'h1de6:    begin Red = 8'h1a;    Green = 8'h1d;    Blue = 8'h3c;
end 13'h1de7:    begin Red = 8'h0b;    Green = 8'h16;    Blue = 8'h34;
end 13'h1de8:    begin Red = 8'h1b;    Green = 8'h20;    Blue = 8'h1c;
end 13'h1de9:    begin Red = 8'h78;    Green = 8'h80;    Blue = 8'h73;
end 13'h1dea:    begin Red = 8'h9f;    Green = 8'h9b;    Blue = 8'h96;
end 13'h1deb:    begin Red = 8'hac;    Green = 8'hf7;    Blue = 8'hfd;
end 13'h1dec:    begin Red = 8'h00;    Green = 8'h00;    Blue = 8'h20;
end 13'h1ded:    begin Red = 8'h34;    Green = 8'h32;    Blue = 8'h1b;
end 13'h1dee:    begin Red = 8'h3a;    Green = 8'h2b;    Blue = 8'h18;
end 13'h1def:    begin Red = 8'h35;    Green = 8'h31;    Blue = 8'h16;
end 13'h1df0:    begin Red = 8'h29;    Green = 8'h22;    Blue = 8'h1c;
end 13'h1df1:    begin Red = 8'h2a;    Green = 8'h26;    Blue = 8'h1b;
end 13'h1df2:    begin Red = 8'h34;    Green = 8'h31;    Blue = 8'h12;
end 13'h1df3:    begin Red = 8'h3c;    Green = 8'h34;    Blue = 8'h1d;
end 13'h1df4:    begin Red = 8'h29;    Green = 8'h15;    Blue = 8'h17;
end 13'h1df5:    begin Red = 8'hc4;    Green = 8'hf9;    Blue = 8'hfd;
end 13'h1df6:    begin Red = 8'ha0;    Green = 8'hff;    Blue = 8'hfe;
end 13'h1df7:    begin Red = 8'h71;    Green = 8'h72;    Blue = 8'h7d;
end 13'h1df8:    begin Red = 8'h70;    Green = 8'h6c;    Blue = 8'h67;
end 13'h1df9:    begin Red = 8'he9;    Green = 8'hdd;    Blue = 8'hb1;
end 13'h1dfa:    begin Red = 8'hea;    Green = 8'hde;    Blue = 8'hbb;
end 13'h1dfb:    begin Red = 8'hea;    Green = 8'he7;    Blue = 8'hc5;
end 13'h1dfc:    begin Red = 8'h02;    Green = 8'he1;    Blue = 8'ha1;
end 13'h1dfd:    begin Red = 8'h04;    Green = 8'h32;    Blue = 8'hb5;
end 13'h1dfe:    begin Red = 8'h04;    Green = 8'h22;    Blue = 8'h70;
end 13'h1dff:    begin Red = 8'h03;    Green = 8'he2;    Blue = 8'h90;
end 13'h1e00:    begin Red = 8'hfa;    Green = 8'hbf;    Blue = 8'h79;
end 13'h1e01:    begin Red = 8'hae;    Green = 8'h93;    Blue = 8'h5b;
end 13'h1e02:    begin Red = 8'h02;    Green = 8'hb1;    Blue = 8'ha0;
end 13'h1e03:    begin Red = 8'h03;    Green = 8'hf2;    Blue = 8'h73;
end 13'h1e04:    begin Red = 8'h03;    Green = 8'hd2;    Blue = 8'h30;
end 13'h1e05:    begin Red = 8'h03;    Green = 8'h81;    Blue = 8'hd0;
end 13'h1e06:    begin Red = 8'h03;    Green = 8'h62;    Blue = 8'h00;
end 13'h1e07:    begin Red = 8'h9c;    Green = 8'h75;    Blue = 8'h4a;
end 13'h1e08:    begin Red = 8'h98;    Green = 8'h88;    Blue = 8'h72;
end 13'h1e09:    begin Red = 8'h4c;    Green = 8'h35;    Blue = 8'h13;
end 13'h1e0a:    begin Red = 8'h04;    Green = 8'h92;    Blue = 8'h66;
end 13'h1e0b:    begin Red = 8'h3a;    Green = 8'hc0;    Blue = 8'hff;
end 13'h1e0c:    begin Red = 8'h3a;    Green = 8'hb6;    Blue = 8'hfc;
end 13'h1e0d:    begin Red = 8'h3b;    Green = 8'hb7;    Blue = 8'hff;
end 13'h1e0e:    begin Red = 8'h54;    Green = 8'h38;    Blue = 8'h11;
end 13'h1e0f:    begin Red = 8'h3d;    Green = 8'hba;    Blue = 8'hfc;
end 13'h1e10:    begin Red = 8'h3d;    Green = 8'hc5;    Blue = 8'hff;
end 13'h1e11:    begin Red = 8'h50;    Green = 8'h49;    Blue = 8'h2f;
end 13'h1e12:    begin Red = 8'h4d;    Green = 8'h47;    Blue = 8'h27;
end 13'h1e13:    begin Red = 8'h02;    Green = 8'h82;    Blue = 8'h15;
end 13'h1e14:    begin Red = 8'h76;    Green = 8'h62;    Blue = 8'h3d;
end 13'h1e15:    begin Red = 8'h99;    Green = 8'h84;    Blue = 8'h59;
end 13'h1e16:    begin Red = 8'h99;    Green = 8'h83;    Blue = 8'h52;
end 13'h1e17:    begin Red = 8'h9a;    Green = 8'h84;    Blue = 8'h55;
end 13'h1e18:    begin Red = 8'h71;    Green = 8'h55;    Blue = 8'h3d;
end 13'h1e19:    begin Red = 8'h79;    Green = 8'h63;    Blue = 8'h3e;
end 13'h1e1a:    begin Red = 8'h79;    Green = 8'h5c;    Blue = 8'h3c;
end 13'h1e1b:    begin Red = 8'h70;    Green = 8'h59;    Blue = 8'h3a;
end 13'h1e1c:    begin Red = 8'h72;    Green = 8'h5e;    Blue = 8'h3d;
end 13'h1e1d:    begin Red = 8'h82;    Green = 8'h61;    Blue = 8'h40;
end 13'h1e1e:    begin Red = 8'h3b;    Green = 8'h2a;    Blue = 8'h20;
end 13'h1e1f:    begin Red = 8'h89;    Green = 8'h7e;    Blue = 8'h88;
end 13'h1e20:    begin Red = 8'hc9;    Green = 8'hff;    Blue = 8'hfe;
end 13'h1e21:    begin Red = 8'hc7;    Green = 8'hfd;    Blue = 8'hff;
end 13'h1e22:    begin Red = 8'h01;    Green = 8'he1;    Blue = 8'h0d;
end 13'h1e23:    begin Red = 8'h4f;    Green = 8'h4d;    Blue = 8'h50;
end 13'h1e24:    begin Red = 8'h55;    Green = 8'h4a;    Blue = 8'h52;
end 13'h1e25:    begin Red = 8'h01;    Green = 8'hf1;    Blue = 8'h6d;
end 13'h1e26:    begin Red = 8'h00;    Green = 8'h34;    Blue = 8'hde;
end 13'h1e27:    begin Red = 8'h64;    Green = 8'h6c;    Blue = 8'h66;
end 13'h1e28:    begin Red = 8'h93;    Green = 8'h7c;    Blue = 8'h5c;
end 13'h1e29:    begin Red = 8'h91;    Green = 8'h7a;    Blue = 8'h58;
end 13'h1e2a:    begin Red = 8'h7b;    Green = 8'h6b;    Blue = 8'h52;
end 13'h1e2b:    begin Red = 8'h95;    Green = 8'h83;    Blue = 8'h5f;
end 13'h1e2c:    begin Red = 8'h4b;    Green = 8'h3e;    Blue = 8'h2e;
end 13'h1e2d:    begin Red = 8'h49;    Green = 8'h3c;    Blue = 8'h2b;
end 13'h1e2e:    begin Red = 8'h3a;    Green = 8'had;    Blue = 8'hfe;
end 13'h1e2f:    begin Red = 8'h37;    Green = 8'h98;    Blue = 8'he5;
end 13'h1e30:    begin Red = 8'h50;    Green = 8'h37;    Blue = 8'h21;
end 13'h1e31:    begin Red = 8'h47;    Green = 8'h3f;    Blue = 8'h2a;
end 13'h1e32:    begin Red = 8'h33;    Green = 8'hac;    Blue = 8'hfd;
end 13'h1e33:    begin Red = 8'h3a;    Green = 8'h97;    Blue = 8'he4;
end 13'h1e34:    begin Red = 8'h7f;    Green = 8'h6f;    Blue = 8'h4d;
end 13'h1e35:    begin Red = 8'he0;    Green = 8'heb;    Blue = 8'hc4;
end 13'h1e36:    begin Red = 8'h44;    Green = 8'h42;    Blue = 8'h43;
end 13'h1e37:    begin Red = 8'h39;    Green = 8'h2b;    Blue = 8'h22;
end 13'h1e38:    begin Red = 8'h43;    Green = 8'h42;    Blue = 8'h3d;
end 13'h1e39:    begin Red = 8'h1b;    Green = 8'h11;    Blue = 8'h10;
end 13'h1e3a:    begin Red = 8'h89;    Green = 8'h7d;    Blue = 8'h7f;
end 13'h1e3b:    begin Red = 8'hb6;    Green = 8'hff;    Blue = 8'hff;
end 13'h1e3c:    begin Red = 8'ha7;    Green = 8'hff;    Blue = 8'hff;
end 13'h1e3d:    begin Red = 8'h01;    Green = 8'hb1;    Blue = 8'h7c;
end 13'h1e3e:    begin Red = 8'h4b;    Green = 8'h47;    Blue = 8'h46;
end 13'h1e3f:    begin Red = 8'h00;    Green = 8'h03;    Blue = 8'h7a;
end 13'h1e40:    begin Red = 8'h71;    Green = 8'h6d;    Blue = 8'h6b;
end 13'h1e41:    begin Red = 8'h81;    Green = 8'h6f;    Blue = 8'h3f;
end 13'h1e42:    begin Red = 8'h83;    Green = 8'h86;    Blue = 8'h88;
end 13'h1e43:    begin Red = 8'h8b;    Green = 8'h82;    Blue = 8'h80;
end 13'h1e44:    begin Red = 8'he5;    Green = 8'he9;    Blue = 8'hc9;
end 13'h1e45:    begin Red = 8'h89;    Green = 8'h88;    Blue = 8'h87;
end 13'h1e46:    begin Red = 8'h92;    Green = 8'h94;    Blue = 8'h7d;
end 13'h1e47:    begin Red = 8'h7c;    Green = 8'h7e;    Blue = 8'h82;
end 13'h1e48:    begin Red = 8'h7e;    Green = 8'h7e;    Blue = 8'h88;
end 13'h1e49:    begin Red = 8'h82;    Green = 8'h84;    Blue = 8'h72;
end 13'h1e4a:    begin Red = 8'h7c;    Green = 8'h87;    Blue = 8'h7d;
end 13'h1e4b:    begin Red = 8'h83;    Green = 8'h7a;    Blue = 8'h88;
end 13'h1e4c:    begin Red = 8'h85;    Green = 8'h83;    Blue = 8'h7c;
end 13'h1e4d:    begin Red = 8'h85;    Green = 8'h80;    Blue = 8'h80;
end 13'h1e4e:    begin Red = 8'he5;    Green = 8'he6;    Blue = 8'hc7;
end 13'h1e4f:    begin Red = 8'h82;    Green = 8'h81;    Blue = 8'h88;
end 13'h1e50:    begin Red = 8'h81;    Green = 8'h84;    Blue = 8'h91;
end 13'h1e51:    begin Red = 8'h81;    Green = 8'h80;    Blue = 8'h85;
end 13'h1e52:    begin Red = 8'h89;    Green = 8'h85;    Blue = 8'h82;
end 13'h1e53:    begin Red = 8'h7e;    Green = 8'h84;    Blue = 8'h8a;
end 13'h1e54:    begin Red = 8'h8a;    Green = 8'h80;    Blue = 8'h8e;
end 13'h1e55:    begin Red = 8'h84;    Green = 8'h80;    Blue = 8'h8c;
end 13'h1e56:    begin Red = 8'h8c;    Green = 8'h85;    Blue = 8'h89;
end 13'h1e57:    begin Red = 8'h7d;    Green = 8'h83;    Blue = 8'h90;
end 13'h1e58:    begin Red = 8'h90;    Green = 8'h82;    Blue = 8'h88;
end 13'h1e59:    begin Red = 8'h77;    Green = 8'h83;    Blue = 8'h85;
end 13'h1e5a:    begin Red = 8'h82;    Green = 8'h88;    Blue = 8'h76;
end 13'h1e5b:    begin Red = 8'h7b;    Green = 8'h79;    Blue = 8'h84;
end 13'h1e5c:    begin Red = 8'h6b;    Green = 8'h69;    Blue = 8'h76;
end 13'h1e5d:    begin Red = 8'h7a;    Green = 8'h82;    Blue = 8'h7c;
end 13'h1e5e:    begin Red = 8'h7d;    Green = 8'h7d;    Blue = 8'h8c;
end 13'h1e5f:    begin Red = 8'h80;    Green = 8'h80;    Blue = 8'h8a;
end 13'h1e60:    begin Red = 8'hb3;    Green = 8'ha1;    Blue = 8'h61;
end 13'h1e61:    begin Red = 8'hb1;    Green = 8'h9f;    Blue = 8'h5f;
end 13'h1e62:    begin Red = 8'hbb;    Green = 8'ha8;    Blue = 8'h57;
end 13'h1e63:    begin Red = 8'hbb;    Green = 8'ha7;    Blue = 8'h51;
end 13'h1e64:    begin Red = 8'hb2;    Green = 8'ha0;    Blue = 8'h65;
end 13'h1e65:    begin Red = 8'hb7;    Green = 8'ha0;    Blue = 8'h5e;
end 13'h1e66:    begin Red = 8'h8a;    Green = 8'h90;    Blue = 8'h83;
end 13'h1e67:    begin Red = 8'hb3;    Green = 8'h9c;    Blue = 8'h53;
end 13'h1e68:    begin Red = 8'hb6;    Green = 8'ha1;    Blue = 8'h55;
end 13'h1e69:    begin Red = 8'hb5;    Green = 8'ha0;    Blue = 8'h59;
end 13'h1e6a:    begin Red = 8'h82;    Green = 8'h87;    Blue = 8'h85;
end 13'h1e6b:    begin Red = 8'h8a;    Green = 8'h84;    Blue = 8'h93;
end 13'h1e6c:    begin Red = 8'hb3;    Green = 8'h9f;    Blue = 8'h5c;
end 13'h1e6d:    begin Red = 8'h95;    Green = 8'h84;    Blue = 8'h82;
end 13'h1e6e:    begin Red = 8'haf;    Green = 8'ha2;    Blue = 8'h5e;
end 13'h1e6f:    begin Red = 8'hb1;    Green = 8'ha2;    Blue = 8'h63;
end 13'h1e70:    begin Red = 8'h88;    Green = 8'h90;    Blue = 8'h88;
end 13'h1e71:    begin Red = 8'h8a;    Green = 8'h84;    Blue = 8'h8b;
end 13'h1e72:    begin Red = 8'hb7;    Green = 8'ha4;    Blue = 8'h50;
end 13'h1e73:    begin Red = 8'ha5;    Green = 8'h95;    Blue = 8'h4a;
end 13'h1e74:    begin Red = 8'h92;    Green = 8'h90;    Blue = 8'h8a;
end 13'h1e75:    begin Red = 8'had;    Green = 8'ha9;    Blue = 8'h92;
end 13'h1e76:    begin Red = 8'h94;    Green = 8'h8d;    Blue = 8'h8b;
end 13'h1e77:    begin Red = 8'h9d;    Green = 8'h8f;    Blue = 8'h87;
end 13'h1e78:    begin Red = 8'h91;    Green = 8'h8e;    Blue = 8'h8d;
end 13'h1e79:    begin Red = 8'h96;    Green = 8'h8e;    Blue = 8'h8d;
end 13'h1e7a:    begin Red = 8'hcb;    Green = 8'hd2;    Blue = 8'hac;
end 13'h1e7b:    begin Red = 8'h8d;    Green = 8'h84;    Blue = 8'h84;
end 13'h1e7c:    begin Red = 8'h94;    Green = 8'h91;    Blue = 8'h92;
end 13'h1e7d:    begin Red = 8'hd4;    Green = 8'hc8;    Blue = 8'hae;
end 13'h1e7e:    begin Red = 8'hd2;    Green = 8'hc7;    Blue = 8'haa;
end 13'h1e7f:    begin Red = 8'hd0;    Green = 8'hc5;    Blue = 8'ha9;
end 13'h1e80:    begin Red = 8'hcf;    Green = 8'hc4;    Blue = 8'ha5;
end 13'h1e81:    begin Red = 8'hcc;    Green = 8'hc1;    Blue = 8'ha3;
end 13'h1e82:    begin Red = 8'hce;    Green = 8'hc2;    Blue = 8'ha1;
end 13'h1e83:    begin Red = 8'hc7;    Green = 8'hba;    Blue = 8'h9d;
end 13'h1e84:    begin Red = 8'hc0;    Green = 8'hb5;    Blue = 8'h99;
end 13'h1e85:    begin Red = 8'hc3;    Green = 8'hb7;    Blue = 8'h96;
end 13'h1e86:    begin Red = 8'hbe;    Green = 8'hb2;    Blue = 8'h93; end
                default: ;
        endcase*/
			end
	 end
    
endmodule
